magic
tech sky130A
magscale 1 2
timestamp 1716529149
<< viali >>
rect 1508 -842 1666 -808
rect 2144 -842 2302 -808
rect 1154 -986 1312 -952
rect 1568 -986 1726 -952
rect 1056 -1552 1092 -1046
rect 2046 -1090 2204 -1056
rect 2470 -1090 2628 -1056
rect 2690 -1446 2724 -1152
<< metal1 >>
rect 1486 -280 1686 -80
rect 1812 -280 2012 -80
rect 2126 -280 2326 -80
rect 245 -303 327 -297
rect 245 -391 327 -385
rect 257 -606 315 -391
rect 1554 -492 1620 -280
rect 1874 -606 1936 -280
rect 2190 -492 2256 -280
rect 3103 -435 3109 -317
rect 3227 -435 3233 -317
rect 2216 -498 2256 -492
rect 3139 -606 3197 -435
rect 257 -664 1562 -606
rect 1608 -664 2200 -606
rect 2244 -664 3197 -606
rect 510 -808 1770 -782
rect 510 -842 1508 -808
rect 1666 -842 1770 -808
rect 510 -888 1770 -842
rect 510 -1348 607 -888
rect 1044 -952 1832 -936
rect 1044 -986 1154 -952
rect 1312 -986 1568 -952
rect 1726 -986 1832 -952
rect 1044 -996 1832 -986
rect 1044 -1046 1104 -996
rect 1044 -1192 1056 -1046
rect 832 -1396 1056 -1192
rect 510 -1704 607 -1445
rect 1044 -1552 1056 -1396
rect 1092 -1192 1104 -1046
rect 1092 -1394 1210 -1192
rect 1256 -1392 1624 -1150
rect 1874 -1180 1936 -664
rect 2034 -808 2446 -790
rect 2034 -842 2144 -808
rect 2302 -842 2446 -808
rect 2034 -884 2446 -842
rect 2180 -924 2264 -884
rect 2180 -1008 2904 -924
rect 2458 -1040 2640 -1008
rect 2036 -1056 2738 -1040
rect 2036 -1090 2046 -1056
rect 2204 -1090 2470 -1056
rect 2628 -1090 2738 -1056
rect 2036 -1102 2738 -1090
rect 2678 -1152 2738 -1102
rect 1674 -1356 2100 -1180
rect 2154 -1356 2522 -1182
rect 2678 -1192 2690 -1152
rect 2572 -1356 2690 -1192
rect 1092 -1552 1104 -1394
rect 1872 -1456 2158 -1396
rect 1872 -1496 1936 -1456
rect 1044 -1566 1104 -1552
rect 1200 -1702 1266 -1502
rect 1614 -1564 1936 -1496
rect 458 -1904 658 -1704
rect 1130 -1902 1330 -1702
rect 1872 -1706 1936 -1564
rect 2516 -1704 2582 -1398
rect 2678 -1446 2690 -1356
rect 2724 -1192 2738 -1152
rect 2820 -1192 2904 -1008
rect 2724 -1310 3050 -1192
rect 2724 -1356 2865 -1310
rect 2724 -1446 2730 -1356
rect 2678 -1460 2730 -1446
rect 2859 -1473 2865 -1356
rect 3028 -1356 3050 -1310
rect 3028 -1473 3034 -1356
rect 2895 -1704 2997 -1473
rect 1814 -1906 2014 -1706
rect 2448 -1904 2648 -1704
rect 2846 -1904 3046 -1704
<< via1 >>
rect 245 -385 327 -303
rect 3109 -435 3227 -317
rect 510 -1445 607 -1348
rect 2865 -1473 3028 -1310
<< metal2 >>
rect 234 -291 339 -282
rect 234 -405 339 -396
rect 3094 -301 3243 -292
rect 3094 -459 3243 -450
rect 469 -1307 648 -1298
rect 469 -1495 648 -1486
rect 2825 -1504 2834 -1279
rect 3059 -1504 3068 -1279
<< via2 >>
rect 234 -303 339 -291
rect 234 -385 245 -303
rect 245 -385 327 -303
rect 327 -385 339 -303
rect 234 -396 339 -385
rect 3094 -317 3243 -301
rect 3094 -435 3109 -317
rect 3109 -435 3227 -317
rect 3227 -435 3243 -317
rect 3094 -450 3243 -435
rect 469 -1348 648 -1307
rect 469 -1445 510 -1348
rect 510 -1445 607 -1348
rect 607 -1445 648 -1348
rect 469 -1486 648 -1445
rect 2834 -1310 3059 -1279
rect 2834 -1473 2865 -1310
rect 2865 -1473 3028 -1310
rect 3028 -1473 3059 -1310
rect 2834 -1504 3059 -1473
<< metal3 >>
rect 209 -265 365 -259
rect 209 -427 365 -421
rect 3070 -277 3267 -271
rect 3070 -480 3267 -474
rect 426 -1523 432 -1270
rect 685 -1523 691 -1270
rect 2815 -1517 2821 -1266
rect 3072 -1517 3078 -1266
<< via3 >>
rect 209 -291 365 -265
rect 209 -396 234 -291
rect 234 -396 339 -291
rect 339 -396 365 -291
rect 209 -421 365 -396
rect 3070 -301 3267 -277
rect 3070 -450 3094 -301
rect 3094 -450 3243 -301
rect 3243 -450 3267 -301
rect 3070 -474 3267 -450
rect 432 -1307 685 -1270
rect 432 -1486 469 -1307
rect 469 -1486 648 -1307
rect 648 -1486 685 -1307
rect 432 -1523 685 -1486
rect 2821 -1279 3072 -1266
rect 2821 -1504 2834 -1279
rect 2834 -1504 3059 -1279
rect 3059 -1504 3072 -1279
rect 2821 -1517 3072 -1504
<< metal4 >>
rect 208 -265 366 -264
rect 208 -421 209 -265
rect 365 -421 978 -265
rect 2644 -277 3270 -274
rect 208 -422 366 -421
rect 2644 -474 3070 -277
rect 3267 -474 3270 -277
rect 2644 -478 3270 -474
rect 432 -1269 685 -774
rect 2821 -1265 3072 -818
rect 2820 -1266 3073 -1265
rect 431 -1270 686 -1269
rect 431 -1523 432 -1270
rect 685 -1523 686 -1270
rect 2820 -1517 2821 -1266
rect 3072 -1517 3073 -1266
rect 2820 -1518 3073 -1517
rect 431 -1524 686 -1523
use sky130_fd_pr__nfet_01v8_64QSBY  sky130_fd_pr__nfet_01v8_64QSBY_0
timestamp 1716528727
transform 1 0 2125 0 1 -1299
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64Z3AY  sky130_fd_pr__nfet_01v8_64Z3AY_0
timestamp 1716517215
transform 1 0 2223 0 1 -599
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64Z3AY  sky130_fd_pr__nfet_01v8_64Z3AY_1
timestamp 1716517215
transform 1 0 1587 0 1 -599
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_LGAKDL  sky130_fd_pr__pfet_01v8_LGAKDL_0
timestamp 1716517215
transform 1 0 1647 0 1 -1300
box -211 -384 211 384
use sky130_fd_pr__cap_mim_m3_1_B4ULDW  XC1
timestamp 1716517215
transform 0 1 916 -1 0 -488
box -396 -460 396 460
use sky130_fd_pr__cap_mim_m3_1_BEWQ6U  XC2
timestamp 1716517215
transform 0 1 2750 -1 0 -520
box -396 -250 396 250
use sky130_fd_pr__pfet_01v8_LGAKDL  XM1
timestamp 1716517215
transform 1 0 1233 0 1 -1300
box -211 -384 211 384
use sky130_fd_pr__nfet_01v8_64QSBY  XM5
timestamp 1716528727
transform 1 0 2549 0 1 -1299
box -211 -279 211 279
<< labels >>
flabel metal1 2126 -280 2326 -80 0 FreeSans 256 0 0 0 s1
port 3 nsew
flabel metal1 1486 -280 1686 -80 0 FreeSans 256 0 0 0 s0
port 2 nsew
flabel metal1 1812 -280 2012 -80 0 FreeSans 256 0 0 0 out
port 4 nsew
flabel metal1 2448 -1904 2648 -1704 0 FreeSans 256 0 0 0 vcont_n
port 6 nsew
flabel metal1 1130 -1902 1330 -1702 0 FreeSans 256 0 0 0 vcont_p
port 1 nsew
flabel metal1 1814 -1906 2014 -1706 0 FreeSans 256 0 0 0 in
port 5 nsew
flabel metal1 832 -1392 1032 -1192 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 458 -1904 658 -1704 0 FreeSans 256 0 0 0 vss
port 7 nsew
flabel metal1 2846 -1904 3046 -1704 0 FreeSans 256 0 0 0 vss
port 7 nsew
<< end >>
