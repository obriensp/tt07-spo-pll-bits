VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_obriensp_pll
  CLASS BLOCK ;
  FOREIGN tt_um_obriensp_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.650000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.350000 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 99.885 72.835 100.055 73.025 ;
        RECT 90.545 72.585 95.640 72.835 ;
        RECT 98.435 72.665 100.195 72.835 ;
        RECT 97.940 72.620 100.195 72.665 ;
        RECT 97.000 72.585 100.195 72.620 ;
        RECT 90.545 72.155 100.195 72.585 ;
        RECT 90.545 71.925 92.565 72.155 ;
        RECT 91.645 71.905 92.565 71.925 ;
        RECT 95.640 71.985 98.870 72.155 ;
        RECT 95.640 71.940 97.930 71.985 ;
        RECT 100.215 71.965 100.645 72.750 ;
        RECT 95.640 71.905 96.990 71.940 ;
      LAYER nwell ;
        RECT 90.350 70.030 100.850 71.635 ;
        RECT 80.000 67.470 102.950 68.630 ;
        RECT 77.750 63.630 102.950 67.470 ;
        RECT 80.000 61.430 102.950 63.630 ;
      LAYER pwell ;
        RECT 125.495 63.535 126.305 63.675 ;
        RECT 125.305 63.365 126.305 63.535 ;
        RECT 125.495 62.305 126.305 63.365 ;
        RECT 80.000 61.020 102.950 61.380 ;
        RECT 77.750 57.230 102.950 61.020 ;
        RECT 80.000 56.330 102.950 57.230 ;
        RECT 125.495 57.095 126.305 62.295 ;
        RECT 125.305 56.925 126.305 57.095 ;
        RECT 125.495 56.785 126.305 56.925 ;
        RECT 125.495 55.720 126.405 56.755 ;
        RECT 125.305 55.550 126.405 55.720 ;
        RECT 125.495 55.405 126.405 55.550 ;
        RECT 125.580 54.955 126.365 55.385 ;
        RECT 125.495 53.875 126.305 54.935 ;
        RECT 125.305 53.705 126.305 53.875 ;
        RECT 125.495 53.565 126.305 53.705 ;
        RECT 125.495 52.500 126.405 53.535 ;
        RECT 125.305 52.330 126.405 52.500 ;
        RECT 125.495 52.185 126.405 52.330 ;
        RECT 125.495 52.030 126.405 52.175 ;
        RECT 125.305 51.860 126.405 52.030 ;
        RECT 125.495 48.285 126.405 51.860 ;
        RECT 125.495 47.890 126.405 48.035 ;
        RECT 125.305 47.720 126.405 47.890 ;
        RECT 125.495 46.685 126.405 47.720 ;
        RECT 125.335 46.340 125.445 46.460 ;
        RECT 125.495 43.755 126.305 46.195 ;
        RECT 125.305 43.585 126.305 43.755 ;
        RECT 125.495 43.445 126.305 43.585 ;
        RECT 125.495 42.375 126.305 43.435 ;
        RECT 125.305 42.205 126.305 42.375 ;
        RECT 125.495 42.065 126.305 42.205 ;
      LAYER nwell ;
        RECT 126.695 41.870 129.525 63.870 ;
      LAYER pwell ;
        RECT 129.915 63.535 130.725 63.675 ;
        RECT 129.915 63.365 130.915 63.535 ;
        RECT 129.915 62.305 130.725 63.365 ;
        RECT 130.770 61.535 130.880 61.695 ;
        RECT 129.815 60.320 130.725 61.355 ;
        RECT 129.815 60.150 130.915 60.320 ;
        RECT 129.815 60.005 130.725 60.150 ;
        RECT 129.815 59.850 130.725 59.995 ;
        RECT 129.815 59.680 130.915 59.850 ;
        RECT 129.815 56.105 130.725 59.680 ;
        RECT 130.775 55.540 130.885 55.660 ;
        RECT 129.855 54.955 130.640 55.385 ;
        RECT 129.815 53.880 130.725 54.915 ;
        RECT 129.815 53.710 130.915 53.880 ;
        RECT 129.815 53.565 130.725 53.710 ;
        RECT 130.775 53.240 130.885 53.360 ;
        RECT 129.915 51.575 130.725 53.095 ;
        RECT 129.915 51.405 130.915 51.575 ;
        RECT 129.915 51.265 130.725 51.405 ;
        RECT 129.815 50.200 130.725 51.235 ;
        RECT 129.815 50.030 130.915 50.200 ;
        RECT 129.815 49.885 130.725 50.030 ;
        RECT 130.745 49.715 130.915 49.735 ;
        RECT 129.905 49.565 130.915 49.715 ;
        RECT 129.905 48.735 130.725 49.565 ;
        RECT 129.815 47.785 130.725 48.735 ;
        RECT 130.775 47.260 130.885 47.380 ;
        RECT 129.915 43.755 130.725 47.115 ;
        RECT 129.915 43.585 130.915 43.755 ;
        RECT 129.915 43.445 130.725 43.585 ;
        RECT 129.915 42.375 130.725 43.435 ;
        RECT 129.915 42.205 130.915 42.375 ;
        RECT 129.915 42.065 130.725 42.205 ;
      LAYER nwell ;
        RECT 107.760 31.330 116.160 36.230 ;
      LAYER pwell ;
        RECT 107.760 28.480 116.120 31.270 ;
      LAYER li1 ;
        RECT 90.540 72.855 100.660 73.025 ;
        RECT 90.625 70.475 90.885 72.685 ;
        RECT 91.135 72.395 91.305 72.855 ;
        RECT 91.475 72.515 92.470 72.685 ;
        RECT 93.000 72.525 93.170 72.685 ;
        RECT 91.475 72.225 91.645 72.515 ;
        RECT 92.300 72.355 92.470 72.515 ;
        RECT 92.640 72.355 93.170 72.525 ;
        RECT 91.075 72.055 91.645 72.225 ;
        RECT 91.815 72.175 91.990 72.345 ;
        RECT 91.075 71.275 91.245 72.055 ;
        RECT 91.815 72.015 92.230 72.175 ;
        RECT 91.820 72.005 92.230 72.015 ;
        RECT 91.555 71.665 92.010 71.835 ;
        RECT 91.075 71.105 91.725 71.275 ;
        RECT 92.640 71.185 92.810 72.355 ;
        RECT 93.515 72.285 93.690 72.615 ;
        RECT 93.860 72.475 94.190 72.855 ;
        RECT 92.980 72.005 93.220 72.175 ;
        RECT 91.055 70.305 91.385 70.685 ;
        RECT 91.555 70.645 91.725 71.105 ;
        RECT 92.025 70.955 92.810 71.185 ;
        RECT 92.025 70.815 92.355 70.955 ;
        RECT 93.050 70.805 93.220 72.005 ;
        RECT 93.515 71.835 93.685 72.285 ;
        RECT 94.460 72.225 94.705 72.645 ;
        RECT 94.880 72.395 95.050 72.855 ;
        RECT 95.220 72.515 96.820 72.685 ;
        RECT 95.220 72.475 95.575 72.515 ;
        RECT 95.810 72.225 95.980 72.345 ;
        RECT 94.460 72.055 95.980 72.225 ;
        RECT 95.810 72.015 95.980 72.055 ;
        RECT 96.150 72.095 96.480 72.345 ;
        RECT 96.650 72.145 96.820 72.515 ;
        RECT 97.110 72.135 97.400 72.855 ;
        RECT 98.110 72.515 99.185 72.685 ;
        RECT 96.150 72.020 96.465 72.095 ;
        RECT 93.395 71.665 93.685 71.835 ;
        RECT 92.510 70.645 92.840 70.685 ;
        RECT 91.555 70.475 92.840 70.645 ;
        RECT 93.010 70.475 93.220 70.805 ;
        RECT 93.515 70.805 93.685 71.665 ;
        RECT 93.855 71.265 94.145 71.945 ;
        RECT 94.620 71.265 94.950 71.885 ;
        RECT 95.155 71.265 95.400 71.885 ;
        RECT 95.795 71.835 96.125 71.845 ;
        RECT 95.740 71.675 96.125 71.835 ;
        RECT 95.740 71.665 95.910 71.675 ;
        RECT 96.295 71.495 96.465 72.020 ;
        RECT 95.705 71.325 96.465 71.495 ;
        RECT 94.470 70.855 95.535 71.025 ;
        RECT 93.515 70.475 93.700 70.805 ;
        RECT 93.870 70.305 94.220 70.685 ;
        RECT 94.470 70.475 94.640 70.855 ;
        RECT 94.810 70.305 95.140 70.685 ;
        RECT 95.365 70.645 95.535 70.855 ;
        RECT 95.705 70.815 96.035 71.325 ;
        RECT 96.205 70.645 96.375 71.155 ;
        RECT 96.635 70.945 96.935 71.945 ;
        RECT 97.580 71.835 97.940 72.510 ;
        RECT 98.110 72.180 98.280 72.515 ;
        RECT 98.450 72.175 98.790 72.345 ;
        RECT 98.500 72.005 98.790 72.175 ;
        RECT 99.015 72.305 99.185 72.515 ;
        RECT 99.355 72.475 99.685 72.855 ;
        RECT 99.855 72.305 100.025 72.680 ;
        RECT 99.015 72.135 100.025 72.305 ;
        RECT 100.285 72.130 100.575 72.855 ;
        RECT 97.580 71.655 98.120 71.835 ;
        RECT 97.580 71.545 97.940 71.655 ;
        RECT 97.135 71.315 97.940 71.545 ;
        RECT 98.620 71.485 98.790 72.005 ;
        RECT 98.155 71.315 98.790 71.485 ;
        RECT 98.960 71.325 99.395 71.945 ;
        RECT 99.705 71.325 100.050 71.945 ;
        RECT 95.365 70.475 96.375 70.645 ;
        RECT 96.635 70.305 96.965 70.685 ;
        RECT 97.135 70.475 97.485 71.315 ;
        RECT 97.655 70.645 97.825 71.145 ;
        RECT 98.155 70.985 98.325 71.315 ;
        RECT 97.995 70.815 98.325 70.985 ;
        RECT 98.495 70.975 100.025 71.145 ;
        RECT 98.495 70.815 98.665 70.975 ;
        RECT 99.015 70.645 99.185 70.805 ;
        RECT 97.655 70.475 99.185 70.645 ;
        RECT 99.355 70.305 99.685 70.685 ;
        RECT 99.855 70.475 100.025 70.975 ;
        RECT 100.285 70.305 100.575 71.470 ;
        RECT 90.540 70.135 100.660 70.305 ;
        RECT 79.530 68.100 80.020 68.590 ;
        RECT 80.400 68.220 82.110 68.390 ;
        RECT 82.950 68.220 84.660 68.390 ;
        RECT 85.500 68.220 87.210 68.390 ;
        RECT 88.050 68.220 89.760 68.390 ;
        RECT 90.600 68.220 92.310 68.390 ;
        RECT 93.150 68.220 94.860 68.390 ;
        RECT 95.700 68.220 97.410 68.390 ;
        RECT 98.250 68.220 99.960 68.390 ;
        RECT 100.800 68.220 102.510 68.390 ;
        RECT 77.930 67.120 79.830 67.290 ;
        RECT 77.930 63.980 78.100 67.120 ;
        RECT 78.500 64.710 78.670 66.750 ;
        RECT 79.090 64.710 79.260 66.750 ;
        RECT 78.715 64.325 79.045 64.495 ;
        RECT 79.660 63.980 79.830 67.120 ;
        RECT 80.800 65.810 80.970 67.850 ;
        RECT 81.540 65.810 81.710 67.850 ;
        RECT 81.030 65.425 81.480 65.595 ;
        RECT 82.110 65.315 82.280 67.985 ;
        RECT 83.350 65.810 83.520 67.850 ;
        RECT 84.090 65.810 84.260 67.850 ;
        RECT 83.580 65.425 84.030 65.595 ;
        RECT 84.660 65.315 84.830 67.985 ;
        RECT 85.900 65.810 86.070 67.850 ;
        RECT 86.640 65.810 86.810 67.850 ;
        RECT 86.130 65.425 86.580 65.595 ;
        RECT 87.210 65.315 87.380 67.985 ;
        RECT 88.450 65.810 88.620 67.850 ;
        RECT 89.190 65.810 89.360 67.850 ;
        RECT 88.680 65.425 89.130 65.595 ;
        RECT 89.760 65.315 89.930 67.985 ;
        RECT 91.000 65.810 91.170 67.850 ;
        RECT 91.740 65.810 91.910 67.850 ;
        RECT 91.230 65.425 91.680 65.595 ;
        RECT 92.310 65.315 92.480 67.985 ;
        RECT 93.550 65.810 93.720 67.850 ;
        RECT 94.290 65.810 94.460 67.850 ;
        RECT 93.780 65.425 94.230 65.595 ;
        RECT 94.860 65.315 95.030 67.985 ;
        RECT 96.100 65.810 96.270 67.850 ;
        RECT 96.840 65.810 97.010 67.850 ;
        RECT 96.330 65.425 96.780 65.595 ;
        RECT 97.410 65.315 97.580 67.985 ;
        RECT 98.650 65.810 98.820 67.850 ;
        RECT 99.390 65.810 99.560 67.850 ;
        RECT 98.880 65.425 99.330 65.595 ;
        RECT 99.960 65.315 100.130 67.985 ;
        RECT 101.200 65.810 101.370 67.850 ;
        RECT 101.940 65.810 102.110 67.850 ;
        RECT 101.430 65.425 101.880 65.595 ;
        RECT 102.510 65.315 102.680 67.985 ;
        RECT 77.930 63.810 79.830 63.980 ;
        RECT 80.800 62.510 80.970 64.550 ;
        RECT 81.540 62.510 81.710 64.550 ;
        RECT 83.350 62.510 83.520 64.550 ;
        RECT 84.090 62.510 84.260 64.550 ;
        RECT 85.900 62.510 86.070 64.550 ;
        RECT 86.640 62.510 86.810 64.550 ;
        RECT 88.450 62.510 88.620 64.550 ;
        RECT 89.190 62.510 89.360 64.550 ;
        RECT 91.000 62.510 91.170 64.550 ;
        RECT 91.740 62.510 91.910 64.550 ;
        RECT 93.550 62.510 93.720 64.550 ;
        RECT 94.290 62.510 94.460 64.550 ;
        RECT 96.100 62.510 96.270 64.550 ;
        RECT 96.840 62.510 97.010 64.550 ;
        RECT 98.650 62.510 98.820 64.550 ;
        RECT 99.390 62.510 99.560 64.550 ;
        RECT 101.200 62.510 101.370 64.550 ;
        RECT 101.940 62.510 102.110 64.550 ;
        RECT 125.305 63.595 125.475 63.680 ;
        RECT 128.025 63.595 128.195 63.680 ;
        RECT 130.745 63.595 130.915 63.680 ;
        RECT 125.305 63.075 126.765 63.595 ;
        RECT 125.305 62.385 126.225 63.075 ;
        RECT 126.935 62.905 129.285 63.595 ;
        RECT 129.455 63.075 130.915 63.595 ;
        RECT 126.395 62.385 129.825 62.905 ;
        RECT 129.995 62.385 130.915 63.075 ;
        RECT 81.030 62.125 81.480 62.295 ;
        RECT 83.580 62.125 84.030 62.295 ;
        RECT 86.130 62.125 86.580 62.295 ;
        RECT 88.680 62.125 89.130 62.295 ;
        RECT 91.230 62.125 91.680 62.295 ;
        RECT 93.780 62.125 94.230 62.295 ;
        RECT 96.330 62.125 96.780 62.295 ;
        RECT 98.880 62.125 99.330 62.295 ;
        RECT 101.430 62.125 101.880 62.295 ;
        RECT 125.305 62.210 125.475 62.385 ;
        RECT 128.025 62.210 128.195 62.385 ;
        RECT 80.230 61.020 82.280 61.190 ;
        RECT 77.930 60.670 79.830 60.840 ;
        RECT 77.930 57.580 78.100 60.670 ;
        RECT 78.500 58.260 78.670 60.300 ;
        RECT 79.090 58.260 79.260 60.300 ;
        RECT 78.715 57.920 79.045 58.090 ;
        RECT 79.660 57.580 79.830 60.670 ;
        RECT 77.930 57.410 79.830 57.580 ;
        RECT 80.230 58.940 80.400 61.020 ;
        RECT 81.030 60.510 81.480 60.680 ;
        RECT 80.800 59.300 80.970 60.340 ;
        RECT 81.540 59.300 81.710 60.340 ;
        RECT 82.110 58.940 82.280 61.020 ;
        RECT 80.230 58.760 82.280 58.940 ;
        RECT 77.430 56.360 77.920 56.850 ;
        RECT 80.230 56.680 80.400 58.760 ;
        RECT 81.030 58.260 81.480 58.430 ;
        RECT 80.800 57.050 80.970 58.090 ;
        RECT 81.540 57.050 81.710 58.090 ;
        RECT 82.110 56.680 82.280 58.760 ;
        RECT 80.230 56.510 82.280 56.680 ;
        RECT 82.780 61.020 84.830 61.190 ;
        RECT 82.780 58.940 82.950 61.020 ;
        RECT 83.580 60.510 84.030 60.680 ;
        RECT 83.350 59.300 83.520 60.340 ;
        RECT 84.090 59.300 84.260 60.340 ;
        RECT 84.660 58.940 84.830 61.020 ;
        RECT 82.780 58.760 84.830 58.940 ;
        RECT 82.780 56.680 82.950 58.760 ;
        RECT 83.580 58.260 84.030 58.430 ;
        RECT 83.350 57.050 83.520 58.090 ;
        RECT 84.090 57.050 84.260 58.090 ;
        RECT 84.660 56.680 84.830 58.760 ;
        RECT 82.780 56.510 84.830 56.680 ;
        RECT 85.330 61.020 87.380 61.190 ;
        RECT 85.330 58.940 85.500 61.020 ;
        RECT 86.130 60.510 86.580 60.680 ;
        RECT 85.900 59.300 86.070 60.340 ;
        RECT 86.640 59.300 86.810 60.340 ;
        RECT 87.210 58.940 87.380 61.020 ;
        RECT 85.330 58.760 87.380 58.940 ;
        RECT 85.330 56.680 85.500 58.760 ;
        RECT 86.130 58.260 86.580 58.430 ;
        RECT 85.900 57.050 86.070 58.090 ;
        RECT 86.640 57.050 86.810 58.090 ;
        RECT 87.210 56.680 87.380 58.760 ;
        RECT 85.330 56.510 87.380 56.680 ;
        RECT 87.880 61.020 89.930 61.190 ;
        RECT 87.880 58.940 88.050 61.020 ;
        RECT 88.680 60.510 89.130 60.680 ;
        RECT 88.450 59.300 88.620 60.340 ;
        RECT 89.190 59.300 89.360 60.340 ;
        RECT 89.760 58.940 89.930 61.020 ;
        RECT 87.880 58.760 89.930 58.940 ;
        RECT 87.880 56.680 88.050 58.760 ;
        RECT 88.680 58.260 89.130 58.430 ;
        RECT 88.450 57.050 88.620 58.090 ;
        RECT 89.190 57.050 89.360 58.090 ;
        RECT 89.760 56.680 89.930 58.760 ;
        RECT 87.880 56.510 89.930 56.680 ;
        RECT 90.430 61.020 92.480 61.190 ;
        RECT 90.430 58.940 90.600 61.020 ;
        RECT 91.230 60.510 91.680 60.680 ;
        RECT 91.000 59.300 91.170 60.340 ;
        RECT 91.740 59.300 91.910 60.340 ;
        RECT 92.310 58.940 92.480 61.020 ;
        RECT 90.430 58.760 92.480 58.940 ;
        RECT 90.430 56.680 90.600 58.760 ;
        RECT 91.230 58.260 91.680 58.430 ;
        RECT 91.000 57.050 91.170 58.090 ;
        RECT 91.740 57.050 91.910 58.090 ;
        RECT 92.310 56.680 92.480 58.760 ;
        RECT 90.430 56.510 92.480 56.680 ;
        RECT 92.980 61.020 95.030 61.190 ;
        RECT 92.980 58.940 93.150 61.020 ;
        RECT 93.780 60.510 94.230 60.680 ;
        RECT 93.550 59.300 93.720 60.340 ;
        RECT 94.290 59.300 94.460 60.340 ;
        RECT 94.860 58.940 95.030 61.020 ;
        RECT 92.980 58.760 95.030 58.940 ;
        RECT 92.980 56.680 93.150 58.760 ;
        RECT 93.780 58.260 94.230 58.430 ;
        RECT 93.550 57.050 93.720 58.090 ;
        RECT 94.290 57.050 94.460 58.090 ;
        RECT 94.860 56.680 95.030 58.760 ;
        RECT 92.980 56.510 95.030 56.680 ;
        RECT 95.530 61.020 97.580 61.190 ;
        RECT 95.530 58.940 95.700 61.020 ;
        RECT 96.330 60.510 96.780 60.680 ;
        RECT 96.100 59.300 96.270 60.340 ;
        RECT 96.840 59.300 97.010 60.340 ;
        RECT 97.410 58.940 97.580 61.020 ;
        RECT 95.530 58.760 97.580 58.940 ;
        RECT 95.530 56.680 95.700 58.760 ;
        RECT 96.330 58.260 96.780 58.430 ;
        RECT 96.100 57.050 96.270 58.090 ;
        RECT 96.840 57.050 97.010 58.090 ;
        RECT 97.410 56.680 97.580 58.760 ;
        RECT 95.530 56.510 97.580 56.680 ;
        RECT 98.080 61.020 100.130 61.190 ;
        RECT 98.080 58.940 98.250 61.020 ;
        RECT 98.880 60.510 99.330 60.680 ;
        RECT 98.650 59.300 98.820 60.340 ;
        RECT 99.390 59.300 99.560 60.340 ;
        RECT 99.960 58.940 100.130 61.020 ;
        RECT 98.080 58.760 100.130 58.940 ;
        RECT 98.080 56.680 98.250 58.760 ;
        RECT 98.880 58.260 99.330 58.430 ;
        RECT 98.650 57.050 98.820 58.090 ;
        RECT 99.390 57.050 99.560 58.090 ;
        RECT 99.960 56.680 100.130 58.760 ;
        RECT 98.080 56.510 100.130 56.680 ;
        RECT 100.630 61.020 102.680 61.190 ;
        RECT 100.630 58.940 100.800 61.020 ;
        RECT 101.430 60.510 101.880 60.680 ;
        RECT 101.200 59.300 101.370 60.340 ;
        RECT 101.940 59.300 102.110 60.340 ;
        RECT 102.510 58.940 102.680 61.020 ;
        RECT 100.630 58.760 102.680 58.940 ;
        RECT 100.630 56.680 100.800 58.760 ;
        RECT 101.430 58.260 101.880 58.430 ;
        RECT 101.200 57.050 101.370 58.090 ;
        RECT 101.940 57.050 102.110 58.090 ;
        RECT 102.510 56.680 102.680 58.760 ;
        RECT 100.630 56.510 102.680 56.680 ;
        RECT 125.305 58.790 126.020 62.210 ;
        RECT 127.590 61.285 128.195 62.210 ;
        RECT 127.590 60.955 129.335 61.285 ;
        RECT 127.590 60.620 128.195 60.955 ;
        RECT 129.505 60.945 129.755 61.295 ;
        RECT 130.745 61.285 130.915 62.385 ;
        RECT 129.935 61.015 130.915 61.285 ;
        RECT 129.935 60.775 130.575 60.845 ;
        RECT 126.340 60.270 128.195 60.620 ;
        RECT 129.165 60.605 130.575 60.775 ;
        RECT 129.165 60.425 129.335 60.605 ;
        RECT 129.935 60.515 130.575 60.605 ;
        RECT 127.590 59.465 128.195 60.270 ;
        RECT 128.380 60.095 129.335 60.425 ;
        RECT 129.505 60.085 129.755 60.435 ;
        RECT 130.745 60.345 130.915 61.015 ;
        RECT 129.935 60.105 130.915 60.345 ;
        RECT 130.745 59.910 130.915 60.105 ;
        RECT 128.365 59.635 129.375 59.910 ;
        RECT 127.590 59.135 128.995 59.465 ;
        RECT 125.305 58.450 126.850 58.790 ;
        RECT 127.590 58.625 128.195 59.135 ;
        RECT 129.165 58.965 129.375 59.635 ;
        RECT 128.365 58.795 129.375 58.965 ;
        RECT 125.305 56.865 126.020 58.450 ;
        RECT 127.590 58.375 128.995 58.625 ;
        RECT 127.590 56.865 128.195 58.375 ;
        RECT 129.165 58.205 129.375 58.795 ;
        RECT 125.305 56.685 125.475 56.865 ;
        RECT 125.305 56.415 126.285 56.685 ;
        RECT 125.305 55.745 125.475 56.415 ;
        RECT 126.465 56.345 126.715 56.695 ;
        RECT 128.025 56.685 128.195 56.865 ;
        RECT 126.885 56.355 128.195 56.685 ;
        RECT 125.645 56.175 126.285 56.245 ;
        RECT 125.645 56.005 127.055 56.175 ;
        RECT 125.645 55.915 126.285 56.005 ;
        RECT 125.305 55.505 126.285 55.745 ;
        RECT 125.305 55.315 125.475 55.505 ;
        RECT 126.465 55.485 126.715 55.835 ;
        RECT 126.885 55.825 127.055 56.005 ;
        RECT 126.885 55.495 127.840 55.825 ;
        RECT 128.025 55.315 128.195 56.355 ;
        RECT 128.365 57.875 129.375 58.205 ;
        RECT 129.555 58.200 129.755 59.860 ;
        RECT 129.925 59.635 130.915 59.910 ;
        RECT 129.925 59.135 130.575 59.465 ;
        RECT 129.925 58.625 130.105 59.135 ;
        RECT 130.745 58.965 130.915 59.635 ;
        RECT 130.275 58.795 130.915 58.965 ;
        RECT 129.925 58.295 130.575 58.625 ;
        RECT 128.365 57.365 128.535 57.875 ;
        RECT 128.705 57.535 129.385 57.705 ;
        RECT 128.365 57.035 128.895 57.365 ;
        RECT 128.365 56.525 128.535 57.035 ;
        RECT 129.085 56.865 129.385 57.535 ;
        RECT 128.705 56.695 129.385 56.865 ;
        RECT 128.365 56.110 128.915 56.525 ;
        RECT 129.085 56.345 129.385 56.695 ;
        RECT 129.555 56.515 129.755 57.880 ;
        RECT 129.925 57.785 130.105 58.295 ;
        RECT 130.745 58.125 130.915 58.795 ;
        RECT 130.275 57.955 130.915 58.125 ;
        RECT 129.925 57.455 130.575 57.785 ;
        RECT 129.925 56.945 130.105 57.455 ;
        RECT 130.745 57.285 130.915 57.955 ;
        RECT 130.275 57.115 130.915 57.285 ;
        RECT 129.925 56.615 130.575 56.945 ;
        RECT 129.925 56.345 130.105 56.615 ;
        RECT 130.745 56.445 130.915 57.115 ;
        RECT 129.085 55.945 130.105 56.345 ;
        RECT 130.275 56.160 130.915 56.445 ;
        RECT 130.745 55.315 130.915 56.160 ;
        RECT 125.305 55.025 126.200 55.315 ;
        RECT 126.860 55.025 129.360 55.315 ;
        RECT 130.020 55.025 130.915 55.315 ;
        RECT 125.305 54.855 125.475 55.025 ;
        RECT 128.025 54.855 128.195 55.025 ;
        RECT 125.305 54.165 126.225 54.855 ;
        RECT 126.395 54.845 128.195 54.855 ;
        RECT 126.395 54.515 129.335 54.845 ;
        RECT 126.395 54.335 128.195 54.515 ;
        RECT 129.505 54.505 129.755 54.855 ;
        RECT 130.745 54.845 130.915 55.025 ;
        RECT 129.935 54.575 130.915 54.845 ;
        RECT 129.935 54.335 130.575 54.405 ;
        RECT 125.305 53.645 126.765 54.165 ;
        RECT 126.935 53.645 128.195 54.335 ;
        RECT 129.165 54.165 130.575 54.335 ;
        RECT 129.165 53.985 129.335 54.165 ;
        RECT 129.935 54.075 130.575 54.165 ;
        RECT 128.380 53.655 129.335 53.985 ;
        RECT 129.505 53.645 129.755 53.995 ;
        RECT 130.745 53.905 130.915 54.575 ;
        RECT 129.935 53.665 130.915 53.905 ;
        RECT 125.305 53.465 125.475 53.645 ;
        RECT 125.305 53.195 126.285 53.465 ;
        RECT 125.305 52.525 125.475 53.195 ;
        RECT 126.465 53.125 126.715 53.475 ;
        RECT 128.025 53.465 128.195 53.645 ;
        RECT 126.885 53.135 128.195 53.465 ;
        RECT 125.645 52.955 126.285 53.025 ;
        RECT 128.025 53.015 128.195 53.135 ;
        RECT 130.745 53.015 130.915 53.665 ;
        RECT 125.645 52.785 127.055 52.955 ;
        RECT 125.645 52.695 126.285 52.785 ;
        RECT 125.305 52.285 126.285 52.525 ;
        RECT 125.305 52.090 125.475 52.285 ;
        RECT 126.465 52.265 126.715 52.615 ;
        RECT 126.885 52.605 127.055 52.785 ;
        RECT 126.885 52.275 127.840 52.605 ;
        RECT 128.025 52.265 129.805 53.015 ;
        RECT 125.305 51.815 126.295 52.090 ;
        RECT 125.305 51.145 125.475 51.815 ;
        RECT 125.645 51.315 126.295 51.645 ;
        RECT 125.305 50.975 125.945 51.145 ;
        RECT 125.305 50.305 125.475 50.975 ;
        RECT 126.115 50.805 126.295 51.315 ;
        RECT 125.645 50.475 126.295 50.805 ;
        RECT 125.305 50.135 125.945 50.305 ;
        RECT 125.305 49.465 125.475 50.135 ;
        RECT 126.115 49.965 126.295 50.475 ;
        RECT 126.465 50.380 126.665 52.040 ;
        RECT 126.845 51.815 127.855 52.090 ;
        RECT 126.845 51.145 127.055 51.815 ;
        RECT 128.025 51.645 129.285 52.265 ;
        RECT 129.975 52.095 130.915 53.015 ;
        RECT 127.225 51.345 129.285 51.645 ;
        RECT 129.455 51.345 130.915 52.095 ;
        RECT 127.225 51.315 128.195 51.345 ;
        RECT 128.025 51.165 128.195 51.315 ;
        RECT 126.845 50.975 127.855 51.145 ;
        RECT 126.845 50.385 127.055 50.975 ;
        RECT 128.025 50.835 129.335 51.165 ;
        RECT 128.025 50.805 128.195 50.835 ;
        RECT 129.505 50.825 129.755 51.175 ;
        RECT 130.745 51.165 130.915 51.345 ;
        RECT 129.935 50.895 130.915 51.165 ;
        RECT 127.225 50.555 128.195 50.805 ;
        RECT 129.935 50.655 130.575 50.725 ;
        RECT 125.645 49.635 126.295 49.965 ;
        RECT 125.305 49.295 125.945 49.465 ;
        RECT 125.305 48.625 125.475 49.295 ;
        RECT 126.115 49.125 126.295 49.635 ;
        RECT 125.645 48.795 126.295 49.125 ;
        RECT 125.305 48.340 125.945 48.625 ;
        RECT 126.115 48.525 126.295 48.795 ;
        RECT 126.465 48.695 126.665 50.060 ;
        RECT 126.845 50.055 127.855 50.385 ;
        RECT 126.835 49.715 127.515 49.885 ;
        RECT 126.835 49.045 127.135 49.715 ;
        RECT 127.685 49.545 127.855 50.055 ;
        RECT 127.325 49.215 127.855 49.545 ;
        RECT 126.835 48.875 127.515 49.045 ;
        RECT 126.835 48.525 127.135 48.875 ;
        RECT 127.685 48.705 127.855 49.215 ;
        RECT 125.305 47.935 125.475 48.340 ;
        RECT 126.115 48.125 127.135 48.525 ;
        RECT 127.305 48.290 127.855 48.705 ;
        RECT 128.025 49.595 128.195 50.555 ;
        RECT 129.165 50.485 130.575 50.655 ;
        RECT 129.165 50.305 129.335 50.485 ;
        RECT 129.935 50.395 130.575 50.485 ;
        RECT 128.380 49.975 129.335 50.305 ;
        RECT 129.505 49.965 129.755 50.315 ;
        RECT 130.745 50.225 130.915 50.895 ;
        RECT 129.935 49.985 130.915 50.225 ;
        RECT 128.025 49.315 128.865 49.595 ;
        RECT 129.145 49.515 129.755 49.780 ;
        RECT 128.025 48.645 128.195 49.315 ;
        RECT 128.535 48.845 129.255 49.145 ;
        RECT 129.505 49.105 129.755 49.515 ;
        RECT 129.925 49.265 130.475 49.595 ;
        RECT 128.025 48.315 128.915 48.645 ;
        RECT 129.085 48.375 129.255 48.845 ;
        RECT 129.505 48.545 129.755 48.885 ;
        RECT 129.925 48.375 130.115 49.265 ;
        RECT 130.745 48.645 130.915 49.985 ;
        RECT 130.285 48.395 130.915 48.645 ;
        RECT 125.305 47.695 126.285 47.935 ;
        RECT 125.305 47.025 125.475 47.695 ;
        RECT 126.465 47.605 126.715 47.955 ;
        RECT 126.885 47.615 127.840 47.945 ;
        RECT 125.645 47.435 126.285 47.525 ;
        RECT 126.885 47.435 127.055 47.615 ;
        RECT 125.645 47.265 127.055 47.435 ;
        RECT 125.645 47.195 126.285 47.265 ;
        RECT 125.305 46.755 126.285 47.025 ;
        RECT 125.305 46.115 125.475 46.755 ;
        RECT 126.465 46.745 126.715 47.095 ;
        RECT 128.025 47.085 128.195 48.315 ;
        RECT 129.085 48.205 130.115 48.375 ;
        RECT 128.365 47.915 128.915 48.125 ;
        RECT 129.505 48.085 129.835 48.205 ;
        RECT 130.285 47.915 130.575 48.225 ;
        RECT 128.365 47.665 130.575 47.915 ;
        RECT 126.885 47.035 128.195 47.085 ;
        RECT 130.745 47.035 130.915 48.395 ;
        RECT 126.885 46.755 129.805 47.035 ;
        RECT 128.025 46.115 129.805 46.755 ;
        RECT 125.305 44.735 126.245 46.115 ;
        RECT 126.415 45.345 129.805 46.115 ;
        RECT 126.415 44.905 129.285 45.345 ;
        RECT 129.975 45.175 130.915 47.035 ;
        RECT 125.305 43.525 126.765 44.735 ;
        RECT 126.935 43.525 129.285 44.905 ;
        RECT 129.455 43.525 130.915 45.175 ;
        RECT 125.305 43.355 125.475 43.525 ;
        RECT 128.025 43.355 128.195 43.525 ;
        RECT 130.745 43.355 130.915 43.525 ;
        RECT 125.305 42.665 126.225 43.355 ;
        RECT 126.395 42.835 129.825 43.355 ;
        RECT 125.305 42.145 126.765 42.665 ;
        RECT 126.935 42.145 129.285 42.835 ;
        RECT 129.995 42.665 130.915 43.355 ;
        RECT 129.455 42.145 130.915 42.665 ;
        RECT 125.305 42.060 125.475 42.145 ;
        RECT 128.025 42.060 128.195 42.145 ;
        RECT 130.745 42.060 130.915 42.145 ;
        RECT 104.860 38.165 105.860 38.450 ;
        RECT 106.460 36.765 107.460 37.050 ;
        RECT 110.390 35.820 111.340 35.990 ;
        RECT 112.490 35.820 113.440 35.990 ;
        RECT 114.590 35.820 115.540 35.990 ;
        RECT 110.700 35.305 111.030 35.475 ;
        RECT 112.800 35.305 113.130 35.475 ;
        RECT 108.340 34.820 109.290 34.990 ;
        RECT 108.510 32.410 108.680 34.450 ;
        RECT 108.950 32.410 109.120 34.450 ;
        RECT 110.560 34.050 110.730 35.090 ;
        RECT 111.000 34.050 111.170 35.090 ;
        RECT 108.650 32.025 108.980 32.195 ;
        RECT 112.660 32.050 112.830 35.090 ;
        RECT 113.100 32.050 113.270 35.090 ;
        RECT 114.760 32.410 114.930 35.450 ;
        RECT 115.200 32.410 115.370 35.450 ;
        RECT 116.160 34.230 116.445 35.230 ;
        RECT 124.645 34.230 124.930 35.230 ;
        RECT 116.160 33.030 116.445 34.030 ;
        RECT 126.445 33.030 126.730 34.030 ;
        RECT 114.900 32.025 115.230 32.195 ;
        RECT 108.650 30.410 108.980 30.580 ;
        RECT 108.510 29.200 108.680 30.240 ;
        RECT 108.950 29.200 109.120 30.240 ;
        RECT 110.610 29.510 110.780 30.550 ;
        RECT 111.050 29.510 111.220 30.550 ;
        RECT 112.660 29.510 112.830 30.550 ;
        RECT 113.100 29.510 113.270 30.550 ;
        RECT 114.900 30.410 115.230 30.580 ;
        RECT 110.750 29.170 111.080 29.340 ;
        RECT 112.800 29.170 113.130 29.340 ;
        RECT 114.760 29.200 114.930 30.240 ;
        RECT 115.200 29.200 115.370 30.240 ;
        RECT 108.340 28.660 109.290 28.830 ;
        RECT 110.440 28.660 111.390 28.830 ;
        RECT 112.490 28.660 113.440 28.830 ;
        RECT 114.590 28.660 115.540 28.830 ;
        RECT 106.460 28.280 107.460 28.565 ;
        RECT 104.860 21.480 105.860 21.765 ;
      LAYER met1 ;
        RECT 77.350 72.730 100.660 73.180 ;
        RECT 90.540 72.700 100.660 72.730 ;
        RECT 83.550 71.575 83.950 71.680 ;
        RECT 90.620 71.575 90.910 72.235 ;
        RECT 92.000 72.160 92.290 72.205 ;
        RECT 92.920 72.160 93.210 72.205 ;
        RECT 98.440 72.160 98.730 72.205 ;
        RECT 92.000 72.020 98.730 72.160 ;
        RECT 92.000 71.975 92.290 72.020 ;
        RECT 92.920 71.975 93.210 72.020 ;
        RECT 98.440 71.975 98.730 72.020 ;
        RECT 91.495 71.820 91.785 71.865 ;
        RECT 93.335 71.820 93.625 71.865 ;
        RECT 91.495 71.680 93.625 71.820 ;
        RECT 91.495 71.635 91.785 71.680 ;
        RECT 93.335 71.635 93.625 71.680 ;
        RECT 93.765 71.580 94.155 71.870 ;
        RECT 94.540 71.580 94.975 71.880 ;
        RECT 95.120 71.580 95.510 71.880 ;
        RECT 95.680 71.820 95.970 71.865 ;
        RECT 97.520 71.820 97.810 71.865 ;
        RECT 98.900 71.840 99.190 71.895 ;
        RECT 95.680 71.680 97.810 71.820 ;
        RECT 95.680 71.635 95.970 71.680 ;
        RECT 97.520 71.635 97.810 71.680 ;
        RECT 83.550 71.430 90.910 71.575 ;
        RECT 83.550 71.330 83.950 71.430 ;
        RECT 90.620 70.925 90.910 71.430 ;
        RECT 96.600 71.525 96.890 71.540 ;
        RECT 96.600 71.265 96.940 71.525 ;
        RECT 98.840 71.430 99.250 71.840 ;
        RECT 99.820 71.735 100.110 71.895 ;
        RECT 98.900 71.265 99.190 71.430 ;
        RECT 99.745 71.325 100.155 71.735 ;
        RECT 99.820 71.265 100.110 71.325 ;
        RECT 96.600 71.245 96.890 71.265 ;
        RECT 92.415 71.140 92.705 71.185 ;
        RECT 95.645 71.140 95.935 71.185 ;
        RECT 92.415 71.000 95.935 71.140 ;
        RECT 92.415 70.955 92.705 71.000 ;
        RECT 95.645 70.955 95.935 71.000 ;
        RECT 90.540 70.430 100.660 70.460 ;
        RECT 79.450 69.980 100.660 70.430 ;
        RECT 79.470 68.630 80.080 68.650 ;
        RECT 77.700 68.080 102.950 68.630 ;
        RECT 79.450 68.040 80.080 68.080 ;
        RECT 79.450 66.730 79.900 68.040 ;
        RECT 81.550 67.830 82.350 68.080 ;
        RECT 84.100 67.830 84.900 68.080 ;
        RECT 86.650 67.830 87.450 68.080 ;
        RECT 89.200 67.830 90.000 68.080 ;
        RECT 91.750 67.830 92.550 68.080 ;
        RECT 94.300 67.830 95.100 68.080 ;
        RECT 96.850 67.830 97.650 68.080 ;
        RECT 99.400 67.830 100.200 68.080 ;
        RECT 101.950 67.830 102.750 68.080 ;
        RECT 78.450 64.530 78.750 66.730 ;
        RECT 79.050 64.730 79.900 66.730 ;
        RECT 78.450 64.080 79.050 64.530 ;
        RECT 79.450 64.230 79.900 64.730 ;
        RECT 80.200 65.830 81.000 67.830 ;
        RECT 81.510 65.830 82.350 67.830 ;
        RECT 82.750 65.830 83.550 67.830 ;
        RECT 84.060 65.830 84.900 67.830 ;
        RECT 85.300 65.830 86.100 67.830 ;
        RECT 86.610 65.830 87.450 67.830 ;
        RECT 87.850 65.830 88.650 67.830 ;
        RECT 89.160 65.830 90.000 67.830 ;
        RECT 90.400 65.830 91.200 67.830 ;
        RECT 91.710 65.830 92.550 67.830 ;
        RECT 92.950 65.830 93.750 67.830 ;
        RECT 94.260 65.830 95.100 67.830 ;
        RECT 95.500 65.830 96.300 67.830 ;
        RECT 96.810 65.830 97.650 67.830 ;
        RECT 98.050 65.830 98.850 67.830 ;
        RECT 99.360 65.830 100.200 67.830 ;
        RECT 100.600 65.830 101.400 67.830 ;
        RECT 101.910 65.830 102.750 67.830 ;
        RECT 117.350 66.400 118.950 66.450 ;
        RECT 80.200 64.530 80.600 65.830 ;
        RECT 80.750 65.130 81.750 65.680 ;
        RECT 82.750 64.530 83.150 65.830 ;
        RECT 83.300 65.130 84.300 65.680 ;
        RECT 85.300 64.530 85.700 65.830 ;
        RECT 85.850 65.130 86.850 65.680 ;
        RECT 87.850 64.530 88.250 65.830 ;
        RECT 88.400 65.130 89.400 65.680 ;
        RECT 90.400 64.530 90.800 65.830 ;
        RECT 90.950 65.130 91.950 65.680 ;
        RECT 92.950 64.530 93.350 65.830 ;
        RECT 93.500 65.130 94.500 65.680 ;
        RECT 95.500 64.530 95.900 65.830 ;
        RECT 96.050 65.130 97.050 65.680 ;
        RECT 98.050 64.530 98.450 65.830 ;
        RECT 98.600 65.130 99.600 65.680 ;
        RECT 100.600 64.530 101.000 65.830 ;
        RECT 101.150 65.130 102.150 65.680 ;
        RECT 117.350 64.900 129.200 66.400 ;
        RECT 117.350 64.850 118.950 64.900 ;
        RECT 78.450 63.230 78.750 64.080 ;
        RECT 78.300 62.730 78.900 63.230 ;
        RECT 78.450 58.330 78.750 62.730 ;
        RECT 80.200 62.530 81.000 64.530 ;
        RECT 81.510 62.530 82.300 64.530 ;
        RECT 82.750 62.530 83.550 64.530 ;
        RECT 84.060 62.530 84.850 64.530 ;
        RECT 85.300 62.530 86.100 64.530 ;
        RECT 86.610 62.530 87.400 64.530 ;
        RECT 87.850 62.530 88.650 64.530 ;
        RECT 89.160 62.530 89.950 64.530 ;
        RECT 90.400 62.530 91.200 64.530 ;
        RECT 91.710 62.530 92.500 64.530 ;
        RECT 92.950 62.530 93.750 64.530 ;
        RECT 94.260 62.530 95.050 64.530 ;
        RECT 95.500 62.530 96.300 64.530 ;
        RECT 96.810 62.530 97.600 64.530 ;
        RECT 98.050 62.530 98.850 64.530 ;
        RECT 99.360 62.530 100.150 64.530 ;
        RECT 100.600 62.530 101.400 64.530 ;
        RECT 101.910 62.530 102.700 64.530 ;
        RECT 81.000 61.680 81.500 62.330 ;
        RECT 80.000 61.130 81.500 61.680 ;
        RECT 81.000 60.480 81.500 61.130 ;
        RECT 81.800 61.680 82.300 62.530 ;
        RECT 83.550 61.680 84.050 62.330 ;
        RECT 81.800 61.130 84.050 61.680 ;
        RECT 79.060 60.230 79.290 60.280 ;
        RECT 79.550 60.230 79.900 60.430 ;
        RECT 81.800 60.330 82.300 61.130 ;
        RECT 83.550 60.480 84.050 61.130 ;
        RECT 84.350 61.680 84.850 62.530 ;
        RECT 86.100 61.680 86.600 62.330 ;
        RECT 86.900 61.680 87.400 62.530 ;
        RECT 88.650 61.680 89.150 62.330 ;
        RECT 84.350 61.130 86.600 61.680 ;
        RECT 86.850 61.130 89.150 61.680 ;
        RECT 84.350 60.330 84.850 61.130 ;
        RECT 86.100 60.480 86.600 61.130 ;
        RECT 86.900 60.330 87.400 61.130 ;
        RECT 88.650 60.480 89.150 61.130 ;
        RECT 89.450 61.680 89.950 62.530 ;
        RECT 91.200 61.680 91.700 62.330 ;
        RECT 92.000 61.680 92.500 62.530 ;
        RECT 93.750 61.680 94.250 62.330 ;
        RECT 89.450 61.130 91.700 61.680 ;
        RECT 91.950 61.130 94.250 61.680 ;
        RECT 89.450 60.330 89.950 61.130 ;
        RECT 91.200 60.480 91.700 61.130 ;
        RECT 92.000 60.330 92.500 61.130 ;
        RECT 93.750 60.480 94.250 61.130 ;
        RECT 94.550 61.680 95.050 62.530 ;
        RECT 96.300 61.680 96.800 62.330 ;
        RECT 97.100 61.680 97.600 62.530 ;
        RECT 98.850 61.680 99.350 62.330 ;
        RECT 94.550 61.130 96.800 61.680 ;
        RECT 97.050 61.130 99.350 61.680 ;
        RECT 94.550 60.330 95.050 61.130 ;
        RECT 96.300 60.480 96.800 61.130 ;
        RECT 97.100 60.330 97.600 61.130 ;
        RECT 98.850 60.480 99.350 61.130 ;
        RECT 99.650 61.680 100.150 62.530 ;
        RECT 101.400 61.680 101.900 62.330 ;
        RECT 102.200 61.680 102.700 62.530 ;
        RECT 99.650 61.130 101.900 61.680 ;
        RECT 102.150 61.130 103.000 61.680 ;
        RECT 99.650 60.330 100.150 61.130 ;
        RECT 101.400 60.480 101.900 61.130 ;
        RECT 102.200 60.330 102.700 61.130 ;
        RECT 79.050 58.330 79.900 60.230 ;
        RECT 78.470 58.280 78.700 58.330 ;
        RECT 79.060 58.280 79.290 58.330 ;
        RECT 78.600 57.680 79.150 58.130 ;
        RECT 77.370 56.880 77.980 56.910 ;
        RECT 79.550 56.880 79.900 58.330 ;
        RECT 80.200 60.320 80.950 60.330 ;
        RECT 81.550 60.320 82.300 60.330 ;
        RECT 80.200 59.330 81.000 60.320 ;
        RECT 80.200 58.080 80.600 59.330 ;
        RECT 80.770 59.320 81.000 59.330 ;
        RECT 81.510 59.330 82.300 60.320 ;
        RECT 82.750 60.320 83.500 60.330 ;
        RECT 84.100 60.320 84.850 60.330 ;
        RECT 82.750 59.330 83.550 60.320 ;
        RECT 81.510 59.320 81.740 59.330 ;
        RECT 80.750 58.230 81.750 58.780 ;
        RECT 82.050 58.080 82.350 58.330 ;
        RECT 80.200 58.070 80.950 58.080 ;
        RECT 81.550 58.070 82.350 58.080 ;
        RECT 80.200 57.080 81.000 58.070 ;
        RECT 80.770 57.070 81.000 57.080 ;
        RECT 81.510 57.070 82.350 58.070 ;
        RECT 82.750 58.080 83.150 59.330 ;
        RECT 83.320 59.320 83.550 59.330 ;
        RECT 84.060 59.330 84.850 60.320 ;
        RECT 85.300 60.320 86.050 60.330 ;
        RECT 86.650 60.320 87.400 60.330 ;
        RECT 85.300 59.330 86.100 60.320 ;
        RECT 84.060 59.320 84.290 59.330 ;
        RECT 83.300 58.230 84.300 58.780 ;
        RECT 84.600 58.080 84.900 58.330 ;
        RECT 82.750 58.070 83.500 58.080 ;
        RECT 84.100 58.070 84.900 58.080 ;
        RECT 82.750 57.080 83.550 58.070 ;
        RECT 83.320 57.070 83.550 57.080 ;
        RECT 84.060 57.070 84.900 58.070 ;
        RECT 85.300 58.080 85.700 59.330 ;
        RECT 85.870 59.320 86.100 59.330 ;
        RECT 86.610 59.330 87.400 60.320 ;
        RECT 87.850 60.320 88.600 60.330 ;
        RECT 89.200 60.320 89.950 60.330 ;
        RECT 87.850 59.330 88.650 60.320 ;
        RECT 86.610 59.320 86.840 59.330 ;
        RECT 85.850 58.230 86.850 58.780 ;
        RECT 87.150 58.080 87.450 58.330 ;
        RECT 85.300 58.070 86.050 58.080 ;
        RECT 86.650 58.070 87.450 58.080 ;
        RECT 85.300 57.080 86.100 58.070 ;
        RECT 85.870 57.070 86.100 57.080 ;
        RECT 86.610 57.070 87.450 58.070 ;
        RECT 87.850 58.080 88.250 59.330 ;
        RECT 88.420 59.320 88.650 59.330 ;
        RECT 89.160 59.330 89.950 60.320 ;
        RECT 90.400 60.320 91.150 60.330 ;
        RECT 91.750 60.320 92.500 60.330 ;
        RECT 90.400 59.330 91.200 60.320 ;
        RECT 89.160 59.320 89.390 59.330 ;
        RECT 88.400 58.230 89.400 58.780 ;
        RECT 89.700 58.080 90.000 58.330 ;
        RECT 87.850 58.070 88.600 58.080 ;
        RECT 89.200 58.070 90.000 58.080 ;
        RECT 87.850 57.080 88.650 58.070 ;
        RECT 88.420 57.070 88.650 57.080 ;
        RECT 89.160 57.070 90.000 58.070 ;
        RECT 90.400 58.080 90.800 59.330 ;
        RECT 90.970 59.320 91.200 59.330 ;
        RECT 91.710 59.330 92.500 60.320 ;
        RECT 92.950 60.320 93.700 60.330 ;
        RECT 94.300 60.320 95.050 60.330 ;
        RECT 92.950 59.330 93.750 60.320 ;
        RECT 91.710 59.320 91.940 59.330 ;
        RECT 90.950 58.230 91.950 58.780 ;
        RECT 92.250 58.080 92.550 58.330 ;
        RECT 90.400 58.070 91.150 58.080 ;
        RECT 91.750 58.070 92.550 58.080 ;
        RECT 90.400 57.080 91.200 58.070 ;
        RECT 90.970 57.070 91.200 57.080 ;
        RECT 91.710 57.070 92.550 58.070 ;
        RECT 92.950 58.080 93.350 59.330 ;
        RECT 93.520 59.320 93.750 59.330 ;
        RECT 94.260 59.330 95.050 60.320 ;
        RECT 95.500 60.320 96.250 60.330 ;
        RECT 96.850 60.320 97.600 60.330 ;
        RECT 95.500 59.330 96.300 60.320 ;
        RECT 94.260 59.320 94.490 59.330 ;
        RECT 93.500 58.230 94.500 58.780 ;
        RECT 94.800 58.080 95.100 58.330 ;
        RECT 92.950 58.070 93.700 58.080 ;
        RECT 94.300 58.070 95.100 58.080 ;
        RECT 92.950 57.080 93.750 58.070 ;
        RECT 93.520 57.070 93.750 57.080 ;
        RECT 94.260 57.070 95.100 58.070 ;
        RECT 95.500 58.080 95.900 59.330 ;
        RECT 96.070 59.320 96.300 59.330 ;
        RECT 96.810 59.330 97.600 60.320 ;
        RECT 98.050 60.320 98.800 60.330 ;
        RECT 99.400 60.320 100.150 60.330 ;
        RECT 98.050 59.330 98.850 60.320 ;
        RECT 96.810 59.320 97.040 59.330 ;
        RECT 96.050 58.230 97.050 58.780 ;
        RECT 97.350 58.080 97.650 58.330 ;
        RECT 95.500 58.070 96.250 58.080 ;
        RECT 96.850 58.070 97.650 58.080 ;
        RECT 95.500 57.080 96.300 58.070 ;
        RECT 96.070 57.070 96.300 57.080 ;
        RECT 96.810 57.070 97.650 58.070 ;
        RECT 98.050 58.080 98.450 59.330 ;
        RECT 98.620 59.320 98.850 59.330 ;
        RECT 99.360 59.330 100.150 60.320 ;
        RECT 100.600 60.320 101.350 60.330 ;
        RECT 101.950 60.320 102.700 60.330 ;
        RECT 100.600 59.330 101.400 60.320 ;
        RECT 99.360 59.320 99.590 59.330 ;
        RECT 98.600 58.230 99.600 58.780 ;
        RECT 99.900 58.080 100.200 58.330 ;
        RECT 98.050 58.070 98.800 58.080 ;
        RECT 99.400 58.070 100.200 58.080 ;
        RECT 98.050 57.080 98.850 58.070 ;
        RECT 98.620 57.070 98.850 57.080 ;
        RECT 99.360 57.070 100.200 58.070 ;
        RECT 100.600 58.080 101.000 59.330 ;
        RECT 101.170 59.320 101.400 59.330 ;
        RECT 101.910 59.330 102.700 60.320 ;
        RECT 101.910 59.320 102.140 59.330 ;
        RECT 101.150 58.230 102.150 58.780 ;
        RECT 102.450 58.080 102.750 58.330 ;
        RECT 100.600 58.070 101.350 58.080 ;
        RECT 101.950 58.070 102.750 58.080 ;
        RECT 100.600 57.080 101.400 58.070 ;
        RECT 101.170 57.070 101.400 57.080 ;
        RECT 101.910 57.070 102.750 58.070 ;
        RECT 81.550 56.880 82.350 57.070 ;
        RECT 84.100 56.880 84.900 57.070 ;
        RECT 86.650 56.880 87.450 57.070 ;
        RECT 89.200 56.880 90.000 57.070 ;
        RECT 91.750 56.880 92.550 57.070 ;
        RECT 94.300 56.880 95.100 57.070 ;
        RECT 96.850 56.880 97.650 57.070 ;
        RECT 99.400 56.880 100.200 57.070 ;
        RECT 101.950 56.880 102.750 57.070 ;
        RECT 77.370 56.330 102.950 56.880 ;
        RECT 77.370 56.300 77.980 56.330 ;
        RECT 97.810 37.580 98.810 44.080 ;
        RECT 99.810 37.580 100.810 52.480 ;
        RECT 117.600 44.300 119.200 44.350 ;
        RECT 125.150 44.300 125.630 63.680 ;
        RECT 127.850 63.200 128.400 64.900 ;
        RECT 126.450 56.390 126.710 56.710 ;
        RECT 126.450 55.470 126.710 55.790 ;
        RECT 127.485 55.485 127.715 55.775 ;
        RECT 127.530 55.330 127.670 55.485 ;
        RECT 127.470 55.010 127.730 55.330 ;
        RECT 126.450 53.170 126.710 53.490 ;
        RECT 126.125 52.725 126.355 53.015 ;
        RECT 126.170 52.020 126.310 52.725 ;
        RECT 126.465 52.480 126.695 52.555 ;
        RECT 126.465 52.340 126.990 52.480 ;
        RECT 126.465 52.265 126.695 52.340 ;
        RECT 126.465 52.020 126.695 52.095 ;
        RECT 126.170 51.880 126.695 52.020 ;
        RECT 126.465 51.805 126.695 51.880 ;
        RECT 126.510 51.190 126.650 51.805 ;
        RECT 126.450 50.870 126.710 51.190 ;
        RECT 126.450 49.720 126.710 49.810 ;
        RECT 126.170 49.580 126.710 49.720 ;
        RECT 126.170 46.960 126.310 49.580 ;
        RECT 126.450 49.490 126.710 49.580 ;
        RECT 126.850 49.350 126.990 52.340 ;
        RECT 127.470 49.950 127.730 50.270 ;
        RECT 126.790 49.030 127.050 49.350 ;
        RECT 126.450 47.650 126.710 47.970 ;
        RECT 127.530 47.955 127.670 49.950 ;
        RECT 127.485 47.665 127.715 47.955 ;
        RECT 126.465 46.960 126.695 47.035 ;
        RECT 126.170 46.820 126.695 46.960 ;
        RECT 126.465 46.745 126.695 46.820 ;
        RECT 117.600 42.800 125.630 44.300 ;
        RECT 117.600 42.750 119.200 42.800 ;
        RECT 125.150 42.060 125.630 42.800 ;
        RECT 127.870 42.060 128.350 63.200 ;
        RECT 129.510 60.990 129.770 61.310 ;
        RECT 128.845 60.085 129.075 60.375 ;
        RECT 129.525 60.085 129.755 60.375 ;
        RECT 128.890 58.920 129.030 60.085 ;
        RECT 129.570 59.380 129.710 60.085 ;
        RECT 129.570 59.240 130.050 59.380 ;
        RECT 129.525 58.920 129.755 58.995 ;
        RECT 128.890 58.780 129.755 58.920 ;
        RECT 128.890 56.710 129.030 58.780 ;
        RECT 129.525 58.705 129.755 58.780 ;
        RECT 129.525 56.865 129.755 57.155 ;
        RECT 128.830 56.390 129.090 56.710 ;
        RECT 128.490 55.470 128.750 55.790 ;
        RECT 128.550 53.935 128.690 55.470 ;
        RECT 129.570 55.330 129.710 56.865 ;
        RECT 129.910 56.250 130.050 59.240 ;
        RECT 129.850 55.930 130.110 56.250 ;
        RECT 129.510 55.010 129.770 55.330 ;
        RECT 129.570 54.855 129.710 55.010 ;
        RECT 129.525 54.565 129.755 54.855 ;
        RECT 128.505 53.645 128.735 53.935 ;
        RECT 129.525 53.860 129.755 53.935 ;
        RECT 129.230 53.720 129.755 53.860 ;
        RECT 128.505 49.965 128.735 50.255 ;
        RECT 128.550 49.810 128.690 49.965 ;
        RECT 128.490 49.490 128.750 49.810 ;
        RECT 129.230 47.970 129.370 53.720 ;
        RECT 129.525 53.645 129.755 53.720 ;
        RECT 129.510 50.870 129.770 51.190 ;
        RECT 129.510 49.950 129.770 50.270 ;
        RECT 129.510 49.030 129.770 49.350 ;
        RECT 129.510 48.570 129.770 48.890 ;
        RECT 129.170 47.650 129.430 47.970 ;
        RECT 130.590 42.060 131.070 63.680 ;
        RECT 104.800 38.100 105.915 38.510 ;
        RECT 97.890 26.850 98.730 37.580 ;
        RECT 99.880 35.915 100.745 37.580 ;
        RECT 105.120 35.915 105.545 38.100 ;
        RECT 108.260 37.580 109.260 38.580 ;
        RECT 115.210 37.580 116.210 38.580 ;
        RECT 106.400 36.705 107.520 37.110 ;
        RECT 108.560 37.000 108.965 37.580 ;
        RECT 115.495 36.985 115.925 37.580 ;
        RECT 128.450 37.550 129.550 38.650 ;
        RECT 107.760 35.915 116.160 36.230 ;
        RECT 99.880 35.730 116.160 35.915 ;
        RECT 99.880 35.050 109.310 35.730 ;
        RECT 108.060 34.730 109.310 35.050 ;
        RECT 110.060 35.080 110.260 35.730 ;
        RECT 110.710 35.280 113.160 35.580 ;
        RECT 110.720 35.275 111.010 35.280 ;
        RECT 111.460 35.080 111.660 35.280 ;
        RECT 112.820 35.275 113.110 35.280 ;
        RECT 114.060 35.080 114.960 35.430 ;
        RECT 108.060 32.430 108.710 34.730 ;
        RECT 108.910 32.430 109.560 34.430 ;
        RECT 108.610 30.380 109.010 32.230 ;
        RECT 109.410 31.930 109.560 32.430 ;
        RECT 110.060 33.680 110.760 35.080 ;
        RECT 110.960 34.080 111.660 35.080 ;
        RECT 110.970 34.070 111.200 34.080 ;
        RECT 112.160 33.680 112.860 35.080 ;
        RECT 110.060 32.080 112.860 33.680 ;
        RECT 113.060 32.430 114.960 35.080 ;
        RECT 115.160 32.830 116.610 35.430 ;
        RECT 124.560 34.910 125.010 35.330 ;
        RECT 128.780 34.965 129.135 37.550 ;
        RECT 128.780 34.910 146.235 34.965 ;
        RECT 124.560 34.610 146.235 34.910 ;
        RECT 124.560 34.555 129.135 34.610 ;
        RECT 124.560 34.130 125.010 34.555 ;
        RECT 126.310 32.930 126.860 34.130 ;
        RECT 115.160 32.430 116.160 32.830 ;
        RECT 135.410 32.580 140.760 34.130 ;
        RECT 145.880 33.430 146.235 34.610 ;
        RECT 145.760 32.880 146.360 33.430 ;
        RECT 113.060 32.080 114.660 32.430 ;
        RECT 112.630 32.070 112.860 32.080 ;
        RECT 113.070 32.070 113.300 32.080 ;
        RECT 114.910 31.930 115.210 32.230 ;
        RECT 109.410 31.630 109.810 31.930 ;
        RECT 114.860 31.630 115.260 31.930 ;
        RECT 109.410 30.230 109.560 31.630 ;
        RECT 107.760 28.880 108.710 30.230 ;
        RECT 108.910 29.230 109.560 30.230 ;
        RECT 110.060 30.780 112.860 31.230 ;
        RECT 110.060 30.530 110.560 30.780 ;
        RECT 110.060 29.530 110.810 30.530 ;
        RECT 108.920 29.220 109.150 29.230 ;
        RECT 110.060 28.880 110.560 29.530 ;
        RECT 111.010 29.380 111.410 30.530 ;
        RECT 112.160 29.530 112.860 30.780 ;
        RECT 114.860 30.630 115.260 30.930 ;
        RECT 113.060 30.230 114.310 30.530 ;
        RECT 114.910 30.380 115.210 30.630 ;
        RECT 115.560 30.230 116.160 32.430 ;
        RECT 113.060 29.530 114.960 30.230 ;
        RECT 110.760 29.080 113.110 29.380 ;
        RECT 113.710 29.230 114.960 29.530 ;
        RECT 115.160 29.230 116.160 30.230 ;
        RECT 114.730 29.220 114.960 29.230 ;
        RECT 115.170 29.220 115.400 29.230 ;
        RECT 107.760 28.625 116.110 28.880 ;
        RECT 106.400 28.480 116.110 28.625 ;
        RECT 106.400 28.220 109.660 28.480 ;
        RECT 107.760 27.430 109.660 28.220 ;
        RECT 137.410 27.430 139.610 32.580 ;
        RECT 107.760 26.850 139.610 27.430 ;
        RECT 97.890 26.010 139.610 26.850 ;
        RECT 107.760 24.880 139.610 26.010 ;
        RECT 104.750 21.420 105.970 21.825 ;
      LAYER met2 ;
        RECT 126.800 85.500 127.200 85.900 ;
        RECT 77.400 72.680 77.950 73.230 ;
        RECT 85.480 72.735 86.070 73.325 ;
        RECT 83.600 71.280 83.900 71.730 ;
        RECT 79.500 69.930 80.050 70.480 ;
        RECT 85.655 68.835 85.900 72.735 ;
        RECT 87.480 72.640 88.070 73.140 ;
        RECT 87.650 71.865 87.905 72.640 ;
        RECT 126.850 72.155 127.150 85.500 ;
        RECT 129.600 81.500 130.000 81.900 ;
        RECT 129.650 72.305 129.950 81.500 ;
        RECT 93.815 71.865 94.105 71.920 ;
        RECT 87.650 71.610 94.105 71.865 ;
        RECT 93.815 71.530 94.105 71.610 ;
        RECT 94.590 71.530 94.880 71.930 ;
        RECT 95.170 71.530 95.460 71.930 ;
        RECT 94.605 69.345 94.850 71.530 ;
        RECT 95.195 70.110 95.430 71.530 ;
        RECT 96.650 71.235 96.910 71.555 ;
        RECT 98.840 71.430 99.250 71.840 ;
        RECT 99.745 71.325 100.155 71.735 ;
        RECT 95.160 69.720 95.460 70.110 ;
        RECT 94.530 69.045 94.920 69.345 ;
        RECT 96.655 68.835 96.900 71.235 ;
        RECT 79.470 68.040 80.080 68.650 ;
        RECT 85.655 68.590 96.900 68.835 ;
        RECT 78.350 65.130 102.950 65.680 ;
        RECT 78.350 62.680 78.850 65.130 ;
        RECT 117.350 64.850 118.950 66.450 ;
        RECT 79.355 63.425 79.855 63.445 ;
        RECT 79.330 58.680 79.880 63.425 ;
        RECT 80.200 61.080 80.950 61.730 ;
        RECT 86.900 61.080 87.650 61.730 ;
        RECT 92.000 61.080 92.750 61.730 ;
        RECT 97.100 61.080 97.850 61.730 ;
        RECT 102.200 61.080 102.950 61.730 ;
        RECT 80.750 58.680 102.950 58.780 ;
        RECT 77.700 58.330 102.950 58.680 ;
        RECT 78.650 57.630 79.100 58.330 ;
        RECT 80.750 58.230 102.950 58.330 ;
        RECT 77.370 56.300 77.980 56.910 ;
        RECT 117.400 52.750 118.900 64.850 ;
        RECT 125.205 60.910 125.575 62.450 ;
        RECT 128.265 61.220 128.635 61.290 ;
        RECT 129.480 61.220 129.800 61.280 ;
        RECT 128.265 61.080 129.800 61.220 ;
        RECT 128.265 61.010 128.635 61.080 ;
        RECT 129.480 61.020 129.800 61.080 ;
        RECT 130.645 60.910 131.015 62.450 ;
        RECT 126.420 56.620 126.740 56.680 ;
        RECT 128.800 56.620 129.120 56.680 ;
        RECT 126.420 56.480 129.120 56.620 ;
        RECT 126.420 56.420 126.740 56.480 ;
        RECT 128.800 56.420 129.120 56.480 ;
        RECT 129.625 56.220 129.995 56.230 ;
        RECT 129.625 55.960 130.140 56.220 ;
        RECT 129.625 55.950 129.995 55.960 ;
        RECT 126.420 55.700 126.740 55.760 ;
        RECT 128.460 55.700 128.780 55.760 ;
        RECT 126.420 55.560 128.780 55.700 ;
        RECT 126.420 55.500 126.740 55.560 ;
        RECT 128.460 55.500 128.780 55.560 ;
        RECT 127.440 55.240 127.760 55.300 ;
        RECT 129.480 55.240 129.800 55.300 ;
        RECT 127.440 55.100 129.800 55.240 ;
        RECT 127.440 55.040 127.760 55.100 ;
        RECT 129.480 55.040 129.800 55.100 ;
        RECT 126.420 53.400 126.740 53.460 ;
        RECT 126.905 53.400 127.275 53.470 ;
        RECT 126.420 53.260 127.275 53.400 ;
        RECT 126.420 53.200 126.740 53.260 ;
        RECT 126.905 53.190 127.275 53.260 ;
        RECT 99.750 51.400 100.850 52.500 ;
        RECT 117.350 51.150 118.950 52.750 ;
        RECT 126.420 51.100 126.740 51.160 ;
        RECT 129.480 51.100 129.800 51.160 ;
        RECT 126.420 50.960 129.800 51.100 ;
        RECT 126.420 50.900 126.740 50.960 ;
        RECT 129.480 50.900 129.800 50.960 ;
        RECT 127.440 50.180 127.760 50.240 ;
        RECT 129.480 50.180 129.800 50.240 ;
        RECT 127.440 50.040 129.800 50.180 ;
        RECT 127.440 49.980 127.760 50.040 ;
        RECT 129.480 49.980 129.800 50.040 ;
        RECT 126.420 49.720 126.740 49.780 ;
        RECT 128.460 49.720 128.780 49.780 ;
        RECT 126.420 49.580 128.780 49.720 ;
        RECT 126.420 49.520 126.740 49.580 ;
        RECT 128.460 49.520 128.780 49.580 ;
        RECT 126.905 49.320 127.275 49.330 ;
        RECT 126.760 49.260 127.275 49.320 ;
        RECT 129.480 49.260 129.800 49.320 ;
        RECT 126.760 49.120 129.800 49.260 ;
        RECT 126.760 49.060 127.275 49.120 ;
        RECT 129.480 49.060 129.800 49.120 ;
        RECT 126.905 49.050 127.275 49.060 ;
        RECT 129.625 48.860 129.995 48.870 ;
        RECT 129.480 48.600 129.995 48.860 ;
        RECT 129.625 48.590 129.995 48.600 ;
        RECT 126.420 47.880 126.740 47.940 ;
        RECT 129.140 47.880 129.460 47.940 ;
        RECT 126.420 47.740 129.460 47.880 ;
        RECT 126.420 47.680 126.740 47.740 ;
        RECT 129.140 47.680 129.460 47.740 ;
        RECT 97.750 43.000 98.850 44.100 ;
        RECT 117.600 42.750 119.200 44.350 ;
        RECT 108.450 37.650 109.150 38.350 ;
        RECT 115.300 37.800 116.000 38.500 ;
        RECT 128.450 37.550 129.550 38.650 ;
        RECT 106.460 36.715 107.460 37.100 ;
        RECT 108.530 37.030 108.995 37.435 ;
        RECT 111.775 37.075 112.075 37.095 ;
        RECT 108.640 31.480 108.885 37.030 ;
        RECT 111.750 35.245 112.100 37.075 ;
        RECT 115.465 37.015 115.955 37.445 ;
        RECT 111.760 35.230 112.060 35.245 ;
        RECT 109.460 31.880 109.760 31.980 ;
        RECT 114.910 31.880 115.210 31.980 ;
        RECT 109.460 31.680 115.210 31.880 ;
        RECT 109.460 31.580 109.760 31.680 ;
        RECT 114.910 31.580 115.210 31.680 ;
        RECT 108.640 31.110 108.960 31.480 ;
        RECT 108.660 31.080 108.960 31.110 ;
        RECT 114.910 30.895 115.210 30.980 ;
        RECT 115.600 30.895 115.825 37.015 ;
        RECT 126.360 32.880 126.810 34.180 ;
        RECT 135.560 32.680 140.610 34.080 ;
        RECT 145.760 32.880 146.360 33.430 ;
        RECT 114.910 30.670 115.825 30.895 ;
        RECT 114.910 30.580 115.210 30.670 ;
        RECT 111.760 29.290 112.060 29.430 ;
        RECT 104.800 21.830 105.920 21.875 ;
        RECT 111.730 21.830 112.140 29.290 ;
        RECT 104.800 21.420 112.140 21.830 ;
        RECT 104.800 21.370 105.920 21.420 ;
      LAYER met3 ;
        RECT 126.750 85.450 127.250 85.950 ;
        RECT 129.550 81.450 130.050 81.950 ;
        RECT 3.405 80.300 4.895 80.325 ;
        RECT 3.400 78.800 80.050 80.300 ;
        RECT 3.405 78.775 4.895 78.800 ;
        RECT 51.485 76.270 52.975 76.295 ;
        RECT 51.480 74.770 77.950 76.270 ;
        RECT 51.485 74.745 52.975 74.770 ;
        RECT 77.400 73.205 77.950 74.770 ;
        RECT 77.350 72.705 78.000 73.205 ;
        RECT 77.400 56.330 77.950 72.705 ;
        RECT 79.500 70.455 80.050 78.800 ;
        RECT 156.415 77.300 157.305 77.325 ;
        RECT 81.550 76.400 157.310 77.300 ;
        RECT 79.450 69.955 80.100 70.455 ;
        RECT 79.500 68.070 80.050 69.955 ;
        RECT 81.550 63.425 82.100 76.400 ;
        RECT 156.415 76.375 157.305 76.400 ;
        RECT 83.560 75.240 83.940 75.560 ;
        RECT 83.600 73.480 83.900 75.240 ;
        RECT 87.560 75.090 87.940 75.410 ;
        RECT 85.640 74.260 85.960 74.640 ;
        RECT 85.650 73.480 85.950 74.260 ;
        RECT 87.600 73.480 87.900 75.090 ;
        RECT 83.500 72.480 84.050 73.480 ;
        RECT 85.500 72.480 86.050 73.480 ;
        RECT 87.500 72.480 88.050 73.480 ;
        RECT 97.350 72.505 100.125 72.855 ;
        RECT 83.595 71.705 83.920 72.480 ;
        RECT 83.550 71.305 83.950 71.705 ;
        RECT 79.330 62.875 82.100 63.425 ;
        RECT 80.150 61.600 81.000 61.705 ;
        RECT 83.595 61.600 83.920 71.305 ;
        RECT 87.100 69.740 95.485 70.090 ;
        RECT 87.100 61.705 87.450 69.740 ;
        RECT 92.200 69.020 94.900 69.370 ;
        RECT 92.200 61.705 92.550 69.020 ;
        RECT 97.350 61.705 97.700 72.505 ;
        RECT 98.870 69.500 99.220 71.810 ;
        RECT 99.775 71.355 100.125 72.505 ;
        RECT 126.825 72.175 127.175 72.525 ;
        RECT 129.625 72.325 129.975 72.675 ;
        RECT 98.870 69.150 102.800 69.500 ;
        RECT 102.450 61.705 102.800 69.150 ;
        RECT 126.850 64.060 127.150 72.175 ;
        RECT 129.650 64.060 129.950 72.325 ;
        RECT 80.150 61.275 83.920 61.600 ;
        RECT 80.150 61.105 81.000 61.275 ;
        RECT 86.850 61.105 87.700 61.705 ;
        RECT 91.950 61.105 92.800 61.705 ;
        RECT 97.050 61.105 97.900 61.705 ;
        RECT 102.150 61.105 103.000 61.705 ;
        RECT 125.225 60.890 125.555 62.470 ;
        RECT 126.790 60.060 127.390 64.060 ;
        RECT 128.285 60.985 128.615 61.315 ;
        RECT 128.300 60.190 128.600 60.985 ;
        RECT 126.940 53.495 127.240 60.060 ;
        RECT 128.290 59.810 128.610 60.190 ;
        RECT 129.510 60.060 130.110 64.060 ;
        RECT 130.665 60.890 130.995 62.470 ;
        RECT 129.650 59.810 129.970 60.060 ;
        RECT 129.645 55.925 129.975 56.255 ;
        RECT 126.925 53.165 127.255 53.495 ;
        RECT 4.405 52.700 5.895 52.725 ;
        RECT 4.400 51.200 118.900 52.700 ;
        RECT 4.405 51.175 5.895 51.200 ;
        RECT 126.925 49.025 127.255 49.355 ;
        RECT 126.940 46.060 127.240 49.025 ;
        RECT 129.660 48.895 129.960 55.925 ;
        RECT 129.645 48.565 129.975 48.895 ;
        RECT 129.660 46.060 129.960 48.565 ;
        RECT 52.505 44.300 53.995 44.325 ;
        RECT 52.500 42.800 119.150 44.300 ;
        RECT 52.505 42.775 53.995 42.800 ;
        RECT 126.790 41.700 127.390 46.060 ;
        RECT 108.500 41.100 127.390 41.700 ;
        RECT 108.500 37.700 109.100 41.100 ;
        RECT 129.510 40.400 130.110 46.060 ;
        RECT 115.350 39.800 130.110 40.400 ;
        RECT 115.350 37.850 115.950 39.800 ;
        RECT 128.555 38.600 129.445 38.625 ;
        RECT 128.550 37.700 129.450 38.600 ;
        RECT 128.555 37.675 129.445 37.700 ;
        RECT 106.410 36.740 112.100 37.075 ;
        RECT 107.310 36.725 112.100 36.740 ;
        RECT 126.310 32.905 126.860 34.155 ;
        RECT 135.510 32.705 140.660 34.055 ;
        RECT 145.760 32.880 146.360 33.430 ;
        RECT 116.210 21.680 138.070 32.080 ;
        RECT 139.660 21.680 151.520 32.080 ;
      LAYER met4 ;
        RECT 3.990 224.400 4.290 224.760 ;
        RECT 7.670 224.400 7.970 224.760 ;
        RECT 11.350 224.400 11.650 224.760 ;
        RECT 15.030 224.400 15.330 224.760 ;
        RECT 18.710 224.400 19.010 224.760 ;
        RECT 22.390 224.400 22.690 224.760 ;
        RECT 26.070 224.400 26.370 224.760 ;
        RECT 29.750 224.400 30.050 224.760 ;
        RECT 33.430 224.400 33.730 224.760 ;
        RECT 37.110 224.400 37.410 224.760 ;
        RECT 40.790 224.400 41.090 224.760 ;
        RECT 44.470 224.400 44.770 224.760 ;
        RECT 48.150 224.400 48.450 224.760 ;
        RECT 51.830 224.400 52.130 224.760 ;
        RECT 55.510 224.400 55.810 224.760 ;
        RECT 59.190 224.400 59.490 224.760 ;
        RECT 62.870 224.400 63.170 224.760 ;
        RECT 66.550 224.400 66.850 224.760 ;
        RECT 70.230 224.400 70.530 224.760 ;
        RECT 73.910 224.400 74.210 224.760 ;
        RECT 77.590 224.400 77.890 224.760 ;
        RECT 81.270 224.400 81.570 224.760 ;
        RECT 84.950 224.400 85.250 224.760 ;
        RECT 2.950 222.850 87.050 224.400 ;
        RECT 88.630 86.250 88.930 224.760 ;
        RECT 83.600 85.950 88.930 86.250 ;
        RECT 2.500 78.800 4.900 80.300 ;
        RECT 50.500 74.770 52.980 76.270 ;
        RECT 83.600 75.565 83.900 85.950 ;
        RECT 126.835 85.850 127.165 85.865 ;
        RECT 136.470 85.850 136.770 224.760 ;
        RECT 126.835 85.550 136.770 85.850 ;
        RECT 126.835 85.535 127.165 85.550 ;
        RECT 129.635 81.850 129.965 81.865 ;
        RECT 140.150 81.850 140.450 224.760 ;
        RECT 129.635 81.550 140.450 81.850 ;
        RECT 129.635 81.535 129.965 81.550 ;
        RECT 143.830 78.550 144.130 224.760 ;
        RECT 87.600 78.250 144.130 78.550 ;
        RECT 83.585 75.235 83.915 75.565 ;
        RECT 87.600 75.415 87.900 78.250 ;
        RECT 87.585 75.085 87.915 75.415 ;
        RECT 85.635 74.600 85.965 74.615 ;
        RECT 147.510 74.600 147.810 224.760 ;
        RECT 85.635 74.300 147.810 74.600 ;
        RECT 85.635 74.285 85.965 74.300 ;
        RECT 125.150 60.880 131.070 62.480 ;
        RECT 128.285 60.150 128.615 60.165 ;
        RECT 129.645 60.150 129.975 60.165 ;
        RECT 128.285 59.850 129.975 60.150 ;
        RECT 128.285 59.835 128.615 59.850 ;
        RECT 129.645 59.835 129.975 59.850 ;
        RECT 2.500 51.200 5.900 52.700 ;
        RECT 50.500 42.800 54.000 44.300 ;
        RECT 128.550 37.700 153.000 38.600 ;
        RECT 126.355 32.925 126.815 34.135 ;
        RECT 126.360 31.685 126.810 32.925 ;
        RECT 135.555 32.740 140.615 34.035 ;
        RECT 145.760 32.880 146.360 33.430 ;
        RECT 135.555 32.725 140.730 32.740 ;
        RECT 137.660 32.020 140.730 32.725 ;
        RECT 116.605 22.075 136.215 31.685 ;
        RECT 137.570 21.840 140.730 32.020 ;
        RECT 145.880 31.685 146.235 32.880 ;
        RECT 141.515 22.075 151.125 31.685 ;
        RECT 137.570 21.830 140.160 21.840 ;
        RECT 137.570 21.740 138.050 21.830 ;
        RECT 139.680 21.740 140.160 21.830 ;
        RECT 152.100 19.250 153.000 37.700 ;
        RECT 134.330 18.350 153.000 19.250 ;
        RECT 134.330 1.000 135.230 18.350 ;
        RECT 156.410 1.000 157.310 77.300 ;
  END
END tt_um_obriensp_pll
END LIBRARY

