magic
tech sky130A
magscale 1 2
timestamp 1717177701
<< viali >>
rect 2789 901 2823 935
rect 1317 833 1351 867
rect 1409 833 1443 867
rect 1593 833 1627 867
rect 1777 833 1811 867
rect 2329 833 2363 867
rect 2513 833 2547 867
rect 2973 833 3007 867
rect 3341 833 3375 867
rect 3617 833 3651 867
rect 3801 833 3835 867
rect 1133 765 1167 799
rect 3617 697 3651 731
rect 1593 629 1627 663
rect 2329 629 2363 663
rect 1133 425 1167 459
rect 2697 425 2731 459
rect 1409 289 1443 323
rect 949 221 983 255
rect 1133 221 1167 255
rect 1501 221 1535 255
rect 1961 221 1995 255
rect 2053 221 2087 255
rect 2237 221 2271 255
rect 2697 221 2731 255
rect 2881 221 2915 255
rect 2145 153 2179 187
<< metal1 >>
rect 0 1114 4324 1136
rect 0 1062 3770 1114
rect 3822 1062 3834 1114
rect 3886 1062 3898 1114
rect 3950 1062 3962 1114
rect 4014 1062 4026 1114
rect 4078 1062 4324 1114
rect 0 1040 4324 1062
rect 2774 892 2780 944
rect 2832 932 2838 944
rect 2832 904 3464 932
rect 2832 892 2838 904
rect 1302 824 1308 876
rect 1360 824 1366 876
rect 1394 824 1400 876
rect 1452 824 1458 876
rect 1578 824 1584 876
rect 1636 824 1642 876
rect 1762 824 1768 876
rect 1820 824 1826 876
rect 2317 867 2375 873
rect 2317 833 2329 867
rect 2363 833 2375 867
rect 2317 827 2375 833
rect 2501 867 2559 873
rect 2501 833 2513 867
rect 2547 864 2559 867
rect 2590 864 2596 876
rect 2547 836 2596 864
rect 2547 833 2559 836
rect 2501 827 2559 833
rect 1118 756 1124 808
rect 1176 796 1182 808
rect 2332 796 2360 827
rect 2590 824 2596 836
rect 2648 864 2654 876
rect 2961 867 3019 873
rect 2961 864 2973 867
rect 2648 836 2973 864
rect 2648 824 2654 836
rect 2961 833 2973 836
rect 3007 833 3019 867
rect 2961 827 3019 833
rect 3329 867 3387 873
rect 3329 833 3341 867
rect 3375 833 3387 867
rect 3436 864 3464 904
rect 3605 867 3663 873
rect 3605 864 3617 867
rect 3436 836 3617 864
rect 3329 827 3387 833
rect 3605 833 3617 836
rect 3651 833 3663 867
rect 3605 827 3663 833
rect 1176 768 2360 796
rect 1176 756 1182 768
rect 2866 688 2872 740
rect 2924 728 2930 740
rect 3344 728 3372 827
rect 3786 824 3792 876
rect 3844 824 3850 876
rect 3605 731 3663 737
rect 3605 728 3617 731
rect 2924 700 3617 728
rect 2924 688 2930 700
rect 3605 697 3617 700
rect 3651 697 3663 731
rect 3605 691 3663 697
rect 1486 620 1492 672
rect 1544 660 1550 672
rect 1581 663 1639 669
rect 1581 660 1593 663
rect 1544 632 1593 660
rect 1544 620 1550 632
rect 1581 629 1593 632
rect 1627 629 1639 663
rect 1581 623 1639 629
rect 2317 663 2375 669
rect 2317 629 2329 663
rect 2363 660 2375 663
rect 2682 660 2688 672
rect 2363 632 2688 660
rect 2363 629 2375 632
rect 2317 623 2375 629
rect 2682 620 2688 632
rect 2740 620 2746 672
rect 0 496 4324 592
rect 1121 459 1179 465
rect 1121 425 1133 459
rect 1167 456 1179 459
rect 1578 456 1584 468
rect 1167 428 1584 456
rect 1167 425 1179 428
rect 1121 419 1179 425
rect 1578 416 1584 428
rect 1636 416 1642 468
rect 2590 416 2596 468
rect 2648 456 2654 468
rect 2685 459 2743 465
rect 2685 456 2697 459
rect 2648 428 2697 456
rect 2648 416 2654 428
rect 2685 425 2697 428
rect 2731 425 2743 459
rect 2685 419 2743 425
rect 1394 280 1400 332
rect 1452 320 1458 332
rect 1452 292 2084 320
rect 1452 280 1458 292
rect 937 255 995 261
rect 937 221 949 255
rect 983 221 995 255
rect 937 215 995 221
rect 952 184 980 215
rect 1118 212 1124 264
rect 1176 212 1182 264
rect 1486 212 1492 264
rect 1544 212 1550 264
rect 1762 212 1768 264
rect 1820 252 1826 264
rect 2056 261 2084 292
rect 1949 255 2007 261
rect 1949 252 1961 255
rect 1820 224 1961 252
rect 1820 212 1826 224
rect 1949 221 1961 224
rect 1995 221 2007 255
rect 1949 215 2007 221
rect 2041 255 2099 261
rect 2041 221 2053 255
rect 2087 221 2099 255
rect 2041 215 2099 221
rect 1504 184 1532 212
rect 952 156 1532 184
rect 1964 184 1992 215
rect 2222 212 2228 264
rect 2280 212 2286 264
rect 2682 212 2688 264
rect 2740 212 2746 264
rect 2866 212 2872 264
rect 2924 212 2930 264
rect 2133 187 2191 193
rect 2133 184 2145 187
rect 1964 156 2145 184
rect 2133 153 2145 156
rect 2179 153 2191 187
rect 2133 147 2191 153
rect 0 26 4324 48
rect 0 -26 3770 26
rect 3822 -26 3834 26
rect 3886 -26 3898 26
rect 3950 -26 3962 26
rect 4014 -26 4026 26
rect 4078 -26 4324 26
rect 0 -48 4324 -26
<< via1 >>
rect 3770 1062 3822 1114
rect 3834 1062 3886 1114
rect 3898 1062 3950 1114
rect 3962 1062 4014 1114
rect 4026 1062 4078 1114
rect 2780 935 2832 944
rect 2780 901 2789 935
rect 2789 901 2823 935
rect 2823 901 2832 935
rect 2780 892 2832 901
rect 1308 867 1360 876
rect 1308 833 1317 867
rect 1317 833 1351 867
rect 1351 833 1360 867
rect 1308 824 1360 833
rect 1400 867 1452 876
rect 1400 833 1409 867
rect 1409 833 1443 867
rect 1443 833 1452 867
rect 1400 824 1452 833
rect 1584 867 1636 876
rect 1584 833 1593 867
rect 1593 833 1627 867
rect 1627 833 1636 867
rect 1584 824 1636 833
rect 1768 867 1820 876
rect 1768 833 1777 867
rect 1777 833 1811 867
rect 1811 833 1820 867
rect 1768 824 1820 833
rect 1124 799 1176 808
rect 1124 765 1133 799
rect 1133 765 1167 799
rect 1167 765 1176 799
rect 2596 824 2648 876
rect 1124 756 1176 765
rect 2872 688 2924 740
rect 3792 867 3844 876
rect 3792 833 3801 867
rect 3801 833 3835 867
rect 3835 833 3844 867
rect 3792 824 3844 833
rect 1492 620 1544 672
rect 2688 620 2740 672
rect 1584 416 1636 468
rect 2596 416 2648 468
rect 1400 323 1452 332
rect 1400 289 1409 323
rect 1409 289 1443 323
rect 1443 289 1452 323
rect 1400 280 1452 289
rect 1124 255 1176 264
rect 1124 221 1133 255
rect 1133 221 1167 255
rect 1167 221 1176 255
rect 1124 212 1176 221
rect 1492 255 1544 264
rect 1492 221 1501 255
rect 1501 221 1535 255
rect 1535 221 1544 255
rect 1492 212 1544 221
rect 1768 212 1820 264
rect 2228 255 2280 264
rect 2228 221 2237 255
rect 2237 221 2271 255
rect 2271 221 2280 255
rect 2228 212 2280 221
rect 2688 255 2740 264
rect 2688 221 2697 255
rect 2697 221 2731 255
rect 2731 221 2740 255
rect 2688 212 2740 221
rect 2872 255 2924 264
rect 2872 221 2881 255
rect 2881 221 2915 255
rect 2915 221 2924 255
rect 2872 212 2924 221
rect 3770 -26 3822 26
rect 3834 -26 3886 26
rect 3898 -26 3950 26
rect 3962 -26 4014 26
rect 4026 -26 4078 26
<< metal2 >>
rect 3770 1116 4078 1125
rect 3770 1114 3776 1116
rect 3832 1114 3856 1116
rect 3912 1114 3936 1116
rect 3992 1114 4016 1116
rect 4072 1114 4078 1116
rect 3832 1062 3834 1114
rect 4014 1062 4016 1114
rect 3770 1060 3776 1062
rect 3832 1060 3856 1062
rect 3912 1060 3936 1062
rect 3992 1060 4016 1062
rect 4072 1060 4078 1062
rect 3770 1051 4078 1060
rect 2780 944 2832 950
rect 1306 912 1362 921
rect 2778 912 2780 921
rect 2832 912 2834 921
rect 1306 847 1308 856
rect 1360 847 1362 856
rect 1400 876 1452 882
rect 1308 818 1360 824
rect 1400 818 1452 824
rect 1584 876 1636 882
rect 1584 818 1636 824
rect 1768 876 1820 882
rect 1768 818 1820 824
rect 2596 876 2648 882
rect 2778 847 2834 856
rect 3792 876 3844 882
rect 2596 818 2648 824
rect 3792 818 3844 824
rect 1124 808 1176 814
rect 1124 750 1176 756
rect 1136 270 1164 750
rect 1412 377 1440 818
rect 1492 672 1544 678
rect 1492 614 1544 620
rect 1398 368 1454 377
rect 1398 303 1400 312
rect 1452 303 1454 312
rect 1400 274 1452 280
rect 1504 270 1532 614
rect 1596 474 1624 818
rect 1584 468 1636 474
rect 1584 410 1636 416
rect 1780 270 1808 818
rect 2608 474 2636 818
rect 2872 740 2924 746
rect 2872 682 2924 688
rect 2688 672 2740 678
rect 2688 614 2740 620
rect 2596 468 2648 474
rect 2596 410 2648 416
rect 2226 368 2282 377
rect 2226 303 2282 312
rect 2240 270 2268 303
rect 2700 270 2728 614
rect 2884 270 2912 682
rect 3804 649 3832 818
rect 3790 640 3846 649
rect 3790 575 3846 584
rect 1124 264 1176 270
rect 1124 206 1176 212
rect 1492 264 1544 270
rect 1492 206 1544 212
rect 1768 264 1820 270
rect 1768 206 1820 212
rect 2228 264 2280 270
rect 2228 206 2280 212
rect 2688 264 2740 270
rect 2688 206 2740 212
rect 2872 264 2924 270
rect 2872 206 2924 212
rect 3770 28 4078 37
rect 3770 26 3776 28
rect 3832 26 3856 28
rect 3912 26 3936 28
rect 3992 26 4016 28
rect 4072 26 4078 28
rect 3832 -26 3834 26
rect 4014 -26 4016 26
rect 3770 -28 3776 -26
rect 3832 -28 3856 -26
rect 3912 -28 3936 -26
rect 3992 -28 4016 -26
rect 4072 -28 4078 -26
rect 3770 -37 4078 -28
<< via2 >>
rect 3776 1114 3832 1116
rect 3856 1114 3912 1116
rect 3936 1114 3992 1116
rect 4016 1114 4072 1116
rect 3776 1062 3822 1114
rect 3822 1062 3832 1114
rect 3856 1062 3886 1114
rect 3886 1062 3898 1114
rect 3898 1062 3912 1114
rect 3936 1062 3950 1114
rect 3950 1062 3962 1114
rect 3962 1062 3992 1114
rect 4016 1062 4026 1114
rect 4026 1062 4072 1114
rect 3776 1060 3832 1062
rect 3856 1060 3912 1062
rect 3936 1060 3992 1062
rect 4016 1060 4072 1062
rect 1306 876 1362 912
rect 2778 892 2780 912
rect 2780 892 2832 912
rect 2832 892 2834 912
rect 1306 856 1308 876
rect 1308 856 1360 876
rect 1360 856 1362 876
rect 2778 856 2834 892
rect 1398 332 1454 368
rect 1398 312 1400 332
rect 1400 312 1452 332
rect 1452 312 1454 332
rect 2226 312 2282 368
rect 3790 584 3846 640
rect 3776 26 3832 28
rect 3856 26 3912 28
rect 3936 26 3992 28
rect 4016 26 4072 28
rect 3776 -26 3822 26
rect 3822 -26 3832 26
rect 3856 -26 3886 26
rect 3886 -26 3898 26
rect 3898 -26 3912 26
rect 3936 -26 3950 26
rect 3950 -26 3962 26
rect 3962 -26 3992 26
rect 4016 -26 4026 26
rect 4026 -26 4072 26
rect 3776 -28 3832 -26
rect 3856 -28 3912 -26
rect 3936 -28 3992 -26
rect 4016 -28 4072 -26
<< metal3 >>
rect 3766 1120 4082 1121
rect 3766 1056 3772 1120
rect 3836 1056 3852 1120
rect 3916 1056 3932 1120
rect 3996 1056 4012 1120
rect 4076 1056 4082 1120
rect 3766 1055 4082 1056
rect 0 914 800 944
rect 1301 914 1367 917
rect 2773 914 2839 917
rect 3600 916 4400 944
rect 0 912 2839 914
rect 0 856 1306 912
rect 1362 856 2778 912
rect 2834 856 2839 912
rect 0 854 2839 856
rect 0 824 800 854
rect 1301 851 1367 854
rect 2773 851 2839 854
rect 3550 852 3556 916
rect 3620 852 4400 916
rect 3600 824 4400 852
rect 3550 580 3556 644
rect 3620 642 3626 644
rect 3785 642 3851 645
rect 3620 640 3851 642
rect 3620 584 3790 640
rect 3846 584 3851 640
rect 3620 582 3851 584
rect 3620 580 3626 582
rect 3785 579 3851 582
rect 0 370 800 400
rect 1393 370 1459 373
rect 0 368 1459 370
rect 0 312 1398 368
rect 1454 312 1459 368
rect 0 310 1459 312
rect 0 280 800 310
rect 1393 307 1459 310
rect 2221 370 2287 373
rect 3600 370 4400 400
rect 2221 368 4400 370
rect 2221 312 2226 368
rect 2282 312 4400 368
rect 2221 310 4400 312
rect 2221 307 2287 310
rect 3600 280 4400 310
rect 3766 32 4082 33
rect 3766 -32 3772 32
rect 3836 -32 3852 32
rect 3916 -32 3932 32
rect 3996 -32 4012 32
rect 4076 -32 4082 32
rect 3766 -33 4082 -32
<< via3 >>
rect 3772 1116 3836 1120
rect 3772 1060 3776 1116
rect 3776 1060 3832 1116
rect 3832 1060 3836 1116
rect 3772 1056 3836 1060
rect 3852 1116 3916 1120
rect 3852 1060 3856 1116
rect 3856 1060 3912 1116
rect 3912 1060 3916 1116
rect 3852 1056 3916 1060
rect 3932 1116 3996 1120
rect 3932 1060 3936 1116
rect 3936 1060 3992 1116
rect 3992 1060 3996 1116
rect 3932 1056 3996 1060
rect 4012 1116 4076 1120
rect 4012 1060 4016 1116
rect 4016 1060 4072 1116
rect 4072 1060 4076 1116
rect 4012 1056 4076 1060
rect 3556 852 3620 916
rect 3556 580 3620 644
rect 3772 28 3836 32
rect 3772 -28 3776 28
rect 3776 -28 3832 28
rect 3832 -28 3836 28
rect 3772 -32 3836 -28
rect 3852 28 3916 32
rect 3852 -28 3856 28
rect 3856 -28 3912 28
rect 3912 -28 3916 28
rect 3852 -32 3916 -28
rect 3932 28 3996 32
rect 3932 -28 3936 28
rect 3936 -28 3992 28
rect 3992 -28 3996 28
rect 3932 -32 3996 -28
rect 4012 28 4076 32
rect 4012 -28 4016 28
rect 4016 -28 4072 28
rect 4072 -28 4076 28
rect 4012 -32 4076 -28
<< metal4 >>
rect 3764 1120 4084 1136
rect 3764 1056 3772 1120
rect 3836 1056 3852 1120
rect 3916 1056 3932 1120
rect 3996 1056 4012 1120
rect 4076 1056 4084 1120
rect 3555 916 3621 917
rect 3555 852 3556 916
rect 3620 852 3621 916
rect 3555 851 3621 852
rect 3558 645 3618 851
rect 3555 644 3621 645
rect 3555 580 3556 644
rect 3620 580 3621 644
rect 3555 579 3621 580
rect 3764 32 4084 1056
rect 3764 -32 3772 32
rect 3836 -32 3852 32
rect 3916 -32 3932 32
rect 3996 -32 4012 32
rect 4076 -32 4084 32
rect 3764 -48 4084 -32
use sky130_fd_sc_hd__and2_1  and0
timestamp 28801
transform -1 0 1564 0 -1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_3
timestamp 28801
transform 1 0 276 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_9
timestamp 28801
transform 1 0 828 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25
timestamp 28801
transform 1 0 2300 0 1 0
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_32
timestamp 1636997256
transform 1 0 2944 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3
timestamp 28801
transform 1 0 276 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_11
timestamp 28801
transform 1 0 1012 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_20
timestamp 28801
transform 1 0 1840 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_24
timestamp 28801
transform 1 0 2208 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_29
timestamp 28801
transform 1 0 2668 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_42
timestamp 28801
transform 1 0 3864 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  l0.n0
timestamp 28801
transform 1 0 2024 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  l0.n1
timestamp 28801
transform -1 0 2024 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  l0.n2
timestamp 28801
transform 1 0 1564 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  l0.n3
timestamp 28801
transform -1 0 1196 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  l1.n0
timestamp 28801
transform 1 0 3588 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  l1.n1
timestamp 28801
transform -1 0 3588 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  l1.n2
timestamp 28801
transform 1 0 2668 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  l1.n3
timestamp 28801
transform 1 0 2300 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_2
timestamp 28801
transform 1 0 0 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 28801
transform -1 0 4324 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_3
timestamp 28801
transform 1 0 0 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 28801
transform -1 0 4324 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_4
timestamp 28801
transform 1 0 2576 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_5
timestamp 28801
transform 1 0 2576 0 -1 1088
box -38 -48 130 592
<< labels >>
flabel metal3 s 3600 824 4400 944 0 FreeSans 480 0 0 0 CLK
port 0 nsew signal input
flabel metal3 s 0 280 800 400 0 FreeSans 480 0 0 0 QA
port 1 nsew signal output
flabel metal3 s 0 824 800 944 0 FreeSans 480 0 0 0 QB
port 2 nsew signal output
flabel metal3 s 3600 280 4400 400 0 FreeSans 480 0 0 0 REF
port 3 nsew signal input
flabel metal4 s 3764 -48 4084 1136 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 -48 28 48 0 FreeSans 224 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 1040 28 1136 0 FreeSans 224 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 496 28 592 0 FreeSans 224 90 0 0 VPWR
port 5 nsew power bidirectional
rlabel metal1 2162 1088 2162 1088 0 VGND
rlabel metal1 2162 544 2162 544 0 VPWR
rlabel metal2 3818 731 3818 731 0 CLK
rlabel via2 1426 323 1426 323 0 QA
rlabel via2 1334 867 1334 867 0 QB
rlabel metal2 2254 289 2254 289 0 REF
rlabel metal1 1748 782 1748 782 0 l0.RESET
rlabel metal1 1978 204 1978 204 0 l0.n0Y
rlabel metal2 1518 442 1518 442 0 l0.n1B
rlabel metal1 1380 442 1380 442 0 l0.n2B
rlabel metal1 3358 782 3358 782 0 l1.n0Y
rlabel metal1 2668 442 2668 442 0 l1.n1B
rlabel metal2 2714 442 2714 442 0 l1.n2B
<< properties >>
string FIXED_BBOX 0 0 4400 1400
<< end >>
