magic
tech sky130A
magscale 1 2
timestamp 1717226440
<< viali >>
rect 5966 -71 6000 -37
rect 5341 -157 5375 -123
rect 5503 -151 5537 -117
rect 6264 -139 6298 -105
rect 6376 -139 6410 -105
rect 6521 -144 6555 -110
rect 7168 -219 7202 19
<< metal1 >>
rect -300 -280 -100 220
rect -300 -390 -260 -280
rect -150 -390 -100 -280
rect -300 -2200 -100 -390
rect 270 180 470 220
rect 270 70 310 180
rect 420 70 470 180
rect 270 -1120 470 70
rect 1010 20 1210 220
rect 1520 20 1720 220
rect 4080 160 4280 220
rect 4080 70 4130 160
rect 4220 70 4280 160
rect 4080 20 4280 70
rect 4610 170 4810 220
rect 4610 80 4670 170
rect 4760 80 4810 170
rect 7216 180 7380 220
rect 5230 124 5233 142
rect 7216 124 7260 180
rect 4610 20 4810 80
rect 7250 70 7260 124
rect 7370 70 7380 180
rect 1055 -410 1145 20
rect 1030 -420 1170 -410
rect 1030 -540 1040 -420
rect 1160 -540 1170 -420
rect 1030 -550 1170 -540
rect 1570 -730 1660 20
rect 7156 19 7214 32
rect 7600 20 7800 220
rect 3434 -20 3566 -14
rect 3434 -140 3440 -20
rect 3560 -58 3566 -20
rect 3560 -102 5372 -58
rect 5940 -80 5950 -20
rect 6010 -25 6020 -20
rect 6010 -80 6022 -25
rect 5944 -83 6022 -80
rect 6242 -93 6320 -92
rect 3560 -140 3566 -102
rect 3434 -146 3566 -140
rect 5319 -111 5372 -102
rect 5319 -123 5397 -111
rect 5481 -117 5559 -105
rect 5481 -122 5503 -117
rect 5319 -157 5341 -123
rect 5375 -157 5397 -123
rect 5319 -169 5397 -157
rect 5461 -151 5503 -122
rect 5537 -151 5559 -117
rect 6236 -149 6246 -93
rect 6298 -149 6320 -93
rect 6242 -151 6320 -149
rect 6354 -94 6432 -93
rect 6354 -105 6378 -94
rect 6354 -139 6376 -105
rect 6354 -150 6378 -139
rect 6430 -150 6440 -94
rect 6500 -98 6510 -90
rect 6499 -150 6510 -98
rect 6570 -150 6580 -90
rect 5461 -163 5559 -151
rect 6354 -152 6432 -150
rect 6499 -156 6577 -150
rect 5461 -211 5498 -163
rect 1854 -248 5498 -211
rect 7156 -219 7168 19
rect 7202 -40 7214 19
rect 7640 -40 7760 20
rect 7202 -160 7760 -40
rect 7202 -219 7214 -160
rect 7156 -231 7214 -219
rect 1854 -414 1927 -248
rect 7250 -324 7260 -280
rect 7230 -390 7260 -324
rect 7370 -390 7380 -280
rect 1830 -420 1950 -414
rect 7230 -420 7380 -390
rect 1830 -546 1950 -540
rect 6219 -555 6225 -485
rect 6295 -555 11090 -485
rect 1570 -735 1960 -730
rect 1570 -845 1845 -735
rect 1955 -845 1961 -735
rect 1570 -850 1960 -845
rect 3300 -1120 3780 -970
rect 7110 -1120 7560 -970
rect 30 -1610 150 -1604
rect 3428 -1608 3572 -1308
rect 1839 -1725 1845 -1615
rect 1955 -1725 1961 -1615
rect 30 -1736 150 -1730
rect 3428 -1752 3952 -1608
rect 7211 -1610 7350 -1311
rect 11020 -1390 11090 -555
rect 5604 -1740 5610 -1620
rect 5730 -1740 5736 -1620
rect 7211 -1749 7740 -1610
rect 9374 -1750 9380 -1630
rect 9500 -1750 9506 -1630
rect -300 -2400 160 -2200
rect 3330 -2400 3780 -2310
rect 7110 -2400 7560 -2310
<< via1 >>
rect -260 -390 -150 -280
rect 310 70 420 180
rect 4130 70 4220 160
rect 4670 80 4760 170
rect 7260 70 7370 180
rect 1040 -540 1160 -420
rect 3440 -140 3560 -20
rect 5950 -37 6010 -20
rect 5950 -71 5966 -37
rect 5966 -71 6000 -37
rect 6000 -71 6010 -37
rect 5950 -80 6010 -71
rect 6246 -105 6298 -93
rect 6246 -139 6264 -105
rect 6264 -139 6298 -105
rect 6246 -149 6298 -139
rect 6378 -105 6430 -94
rect 6378 -139 6410 -105
rect 6410 -139 6430 -105
rect 6378 -150 6430 -139
rect 6510 -110 6570 -90
rect 6510 -144 6521 -110
rect 6521 -144 6555 -110
rect 6555 -144 6570 -110
rect 6510 -150 6570 -144
rect 7260 -390 7370 -280
rect 1830 -540 1950 -420
rect 6225 -555 6295 -485
rect 1845 -845 1955 -735
rect 30 -1730 150 -1610
rect 1845 -1725 1955 -1615
rect 5610 -1740 5730 -1620
rect 9380 -1750 9500 -1630
<< metal2 >>
rect 310 180 420 190
rect 7260 180 7370 190
rect 4670 170 4760 180
rect 310 60 420 70
rect 4130 160 4220 170
rect 4760 147 4770 170
rect 4760 105 6557 147
rect 4760 80 4770 105
rect 4670 70 4760 80
rect 4130 0 4220 70
rect 3434 -20 3566 -14
rect 3434 -140 3440 -20
rect 3560 -140 3566 -20
rect 4135 -28 4205 0
rect 5950 -20 6010 -10
rect 4135 -72 5950 -28
rect 6515 -80 6557 105
rect 7260 60 7370 70
rect 5950 -90 6010 -80
rect 6246 -85 6298 -83
rect 3434 -146 3566 -140
rect 6225 -93 6298 -85
rect -260 -280 -150 -270
rect -260 -400 -150 -390
rect 1030 -420 1170 -410
rect 70 -540 1040 -420
rect 1160 -540 1830 -420
rect 1950 -540 1956 -420
rect 70 -680 190 -540
rect 1030 -550 1170 -540
rect -180 -800 190 -680
rect 1845 -735 1955 -729
rect -180 -1610 -60 -800
rect -180 -1730 30 -1610
rect 150 -1730 156 -1610
rect 1845 -1615 1955 -845
rect 3440 -1330 3560 -146
rect 6225 -149 6246 -93
rect 6378 -94 6430 -84
rect 6225 -159 6298 -149
rect 6375 -150 6378 -95
rect 6510 -90 6570 -80
rect 6430 -150 6445 -95
rect 6225 -485 6295 -159
rect 6225 -561 6295 -555
rect 6375 -830 6445 -150
rect 6510 -160 6570 -150
rect 7260 -280 7370 -270
rect 7260 -400 7370 -390
rect 6375 -900 7310 -830
rect 7240 -1405 7310 -900
rect 1845 -1731 1955 -1725
rect 5610 -1620 5730 -1614
rect 3450 -2500 3570 -1960
rect 5610 -2500 5730 -1740
rect 9380 -1630 9500 -1624
rect 3450 -2620 5730 -2500
rect 7220 -2500 7340 -1960
rect 9380 -2500 9500 -1750
rect 7220 -2620 9500 -2500
<< via2 >>
rect 310 70 420 180
rect 7260 70 7370 180
rect -260 -390 -150 -280
rect 7260 -390 7370 -280
<< metal3 >>
rect 300 180 430 185
rect 7250 180 7380 185
rect 300 70 310 180
rect 420 70 7260 180
rect 7370 70 7380 180
rect 300 65 430 70
rect 7250 65 7380 70
rect -270 -280 -140 -275
rect 7250 -280 7380 -275
rect -270 -390 -260 -280
rect -150 -390 7260 -280
rect 7370 -390 7380 -280
rect -270 -395 -140 -390
rect 7250 -395 7380 -390
use clkdiv2  x4
timestamp 1717213418
transform 1 0 0 0 1 -400
box 0 -2000 3600 -570
use clkdiv2  x5
timestamp 1717213418
transform 1 0 3780 0 1 -400
box 0 -2000 3600 -570
use clkdiv2  x6
timestamp 1717213418
transform 1 0 7560 0 1 -400
box 0 -2000 3600 -570
use sky130_fd_sc_hd__tapvpwrvgnd_1  x8
timestamp 1717194565
transform 1 0 5208 0 1 -372
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  x11
timestamp 1717194565
transform 1 0 5298 0 1 -372
box -38 -48 1970 592
<< labels >>
flabel metal1 1010 20 1210 220 0 FreeSans 256 0 0 0 clk
port 5 nsew
flabel metal1 1520 20 1720 220 0 FreeSans 256 0 0 0 clk_n
port 6 nsew
flabel metal1 -300 20 -100 220 0 FreeSans 256 0 0 0 vss
port 2 nsew
flabel metal1 270 20 470 220 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 7600 20 7800 220 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 4610 20 4810 220 0 FreeSans 256 0 0 0 s1
port 4 nsew
flabel metal1 4080 20 4280 220 0 FreeSans 256 0 0 0 s0
port 3 nsew
<< end >>
