magic
tech sky130A
magscale 1 2
timestamp 1717173898
<< metal3 >>
rect 681 16060 979 16065
rect 680 16059 16010 16060
rect 680 15761 681 16059
rect 979 15761 16010 16059
rect 680 15760 16010 15761
rect 681 15755 979 15760
rect 10297 15254 10595 15259
rect 10296 15253 15590 15254
rect 10296 14955 10297 15253
rect 10595 14955 15590 15253
rect 10296 14954 15590 14955
rect 10297 14949 10595 14954
rect 15480 14670 15590 14954
rect 15900 14650 16010 15760
rect 31283 15460 31461 15465
rect 16310 15459 31462 15460
rect 16310 15281 31283 15459
rect 31461 15281 31462 15459
rect 16310 15280 31462 15281
rect 16310 14510 16420 15280
rect 31283 15275 31461 15280
rect 16712 15048 16718 15112
rect 16782 15048 16788 15112
rect 16720 14580 16780 15048
rect 17512 15018 17518 15082
rect 17582 15018 17588 15082
rect 17128 14922 17192 14928
rect 17128 14852 17192 14858
rect 17130 14570 17190 14852
rect 17520 14590 17580 15018
<< via3 >>
rect 681 15761 979 16059
rect 10297 14955 10595 15253
rect 31283 15281 31461 15459
rect 16718 15048 16782 15112
rect 17518 15018 17582 15082
rect 17128 14858 17192 14922
<< metal4 >>
rect 798 44880 858 45152
rect 1534 44880 1594 45152
rect 2270 44880 2330 45152
rect 3006 44880 3066 45152
rect 3742 44880 3802 45152
rect 4478 44880 4538 45152
rect 5214 44880 5274 45152
rect 5950 44880 6010 45152
rect 6686 44880 6746 45152
rect 7422 44880 7482 45152
rect 8158 44880 8218 45152
rect 8894 44880 8954 45152
rect 9630 44880 9690 45152
rect 10366 44880 10426 45152
rect 11102 44880 11162 45152
rect 11838 44880 11898 45152
rect 12574 44880 12634 45152
rect 13310 44880 13370 45152
rect 14046 44880 14106 45152
rect 14782 44880 14842 45152
rect 15518 44880 15578 45152
rect 16254 44880 16314 45152
rect 16990 44880 17050 45152
rect 590 44570 17410 44880
rect 200 16060 500 44152
rect 200 16059 980 16060
rect 200 15761 681 16059
rect 979 15761 980 16059
rect 200 15760 980 15761
rect 200 1000 500 15760
rect 9800 15254 10100 44152
rect 17726 17250 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 16720 17190 17786 17250
rect 9800 15253 10596 15254
rect 9800 14955 10297 15253
rect 10595 14955 10596 15253
rect 16720 15113 16780 17190
rect 28766 15710 28826 45152
rect 17520 15650 28826 15710
rect 16717 15112 16783 15113
rect 16717 15048 16718 15112
rect 16782 15048 16783 15112
rect 17520 15083 17580 15650
rect 16717 15047 16783 15048
rect 17517 15082 17583 15083
rect 17517 15018 17518 15082
rect 17582 15018 17583 15082
rect 17517 15017 17583 15018
rect 9800 14954 10596 14955
rect 9800 1000 10100 14954
rect 17127 14922 17193 14923
rect 17127 14858 17128 14922
rect 17192 14920 17193 14922
rect 29502 14920 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 17192 14860 29562 14920
rect 31282 15459 31462 15460
rect 31282 15281 31283 15459
rect 31461 15281 31462 15459
rect 17192 14858 17193 14860
rect 17127 14857 17193 14858
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 15281
use vco  vco_0
timestamp 1717119155
transform 1 0 16000 0 1 12466
box -530 -1206 4600 2230
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
