magic
tech sky130A
magscale 1 2
timestamp 1717186736
<< nwell >>
rect 3840 580 5520 1560
<< viali >>
rect 3260 1947 3460 2004
rect 3580 1667 3780 1724
rect 4382 1478 4540 1512
rect 4802 1478 4960 1512
rect 5222 1478 5380 1512
rect 3972 1278 4130 1312
rect 5520 1160 5577 1360
rect 7217 1160 7274 1360
rect 5520 920 5577 1120
rect 7577 920 7634 1120
rect 3972 46 4130 80
rect 4392 46 4550 80
rect 4802 46 4960 80
rect 5222 46 5380 80
rect 3580 -30 3780 27
rect 3260 -1390 3460 -1333
<< metal1 >>
rect 1850 1830 2050 2030
rect 2250 1830 2450 2030
rect 3248 2004 3471 2016
rect 3248 1947 3260 2004
rect 3460 1947 3471 2004
rect 3248 1934 3471 1947
rect 1866 -316 2034 1830
rect 2264 1497 2437 1830
rect 3312 1497 3397 1934
rect 3940 1830 4140 2030
rect 5330 1830 5530 2030
rect 7990 1830 8190 2030
rect 4000 1801 4081 1830
rect 3568 1724 3792 1736
rect 3568 1667 3580 1724
rect 3780 1667 3792 1724
rect 4000 1714 4081 1720
rect 5387 1803 5473 1830
rect 5387 1711 5473 1717
rect 3568 1655 3792 1667
rect 3840 1512 5520 1560
rect 3840 1497 4382 1512
rect 2264 1478 4382 1497
rect 4540 1478 4802 1512
rect 4960 1478 5222 1512
rect 5380 1478 5520 1512
rect 2264 1460 5520 1478
rect 2264 1324 4150 1460
rect 3900 1312 4150 1324
rect 3900 1278 3972 1312
rect 4130 1278 4150 1312
rect 3900 1260 4150 1278
rect 4300 1330 4340 1460
rect 4430 1370 4640 1430
rect 4700 1370 4920 1430
rect 4580 1330 4620 1370
rect 5100 1330 5280 1400
rect 3900 800 4030 1260
rect 4070 800 4200 1200
rect 4010 600 4090 760
rect 4010 540 4020 600
rect 4080 540 4090 600
rect 4010 390 4090 540
rect 4170 700 4200 800
rect 4300 1050 4440 1330
rect 4480 1130 4620 1330
rect 4720 1050 4860 1330
rect 4300 730 4860 1050
rect 4900 800 5280 1330
rect 5320 1360 5610 1400
rect 5320 1160 5520 1360
rect 5577 1160 5610 1360
rect 5320 1120 5610 1160
rect 7200 1360 7290 1380
rect 7200 1160 7217 1360
rect 7274 1296 7290 1360
rect 8044 1307 8115 1830
rect 8044 1296 11535 1307
rect 7274 1236 11535 1296
rect 7274 1225 8115 1236
rect 7274 1160 7290 1225
rect 7200 1140 7290 1160
rect 5320 920 5520 1120
rect 5577 920 5610 1120
rect 5320 880 5610 920
rect 7550 900 7560 1140
rect 7650 900 7660 1140
rect 9370 1120 10440 1140
rect 5320 800 5520 880
rect 9370 860 9400 1120
rect 10410 860 10440 1120
rect 11464 1000 11535 1236
rect 11440 976 11560 1000
rect 11440 905 11464 976
rect 11535 905 11560 976
rect 11440 890 11560 905
rect 9370 830 10440 860
rect 4900 730 5220 800
rect 5270 700 5330 760
rect 4170 640 4180 700
rect 4240 640 4250 700
rect 5260 640 5270 700
rect 5330 640 5340 700
rect 4170 360 4200 640
rect 3840 90 4030 360
rect 4070 160 4200 360
rect 4300 470 4860 560
rect 4300 420 4400 470
rect 4300 220 4450 420
rect 4300 90 4400 220
rect 4490 190 4570 420
rect 4720 220 4860 470
rect 5260 440 5270 500
rect 5330 440 5340 500
rect 4900 360 5150 420
rect 5270 390 5330 440
rect 5400 360 5520 800
rect 4900 220 5280 360
rect 4440 130 4640 190
rect 4700 130 4910 190
rect 5030 160 5280 220
rect 5320 160 5520 360
rect 3840 80 5510 90
rect 3840 46 3972 80
rect 4130 46 4392 80
rect 4550 46 4802 80
rect 4960 46 5222 80
rect 5380 46 5510 80
rect 3840 39 5510 46
rect 3568 27 5510 39
rect 3568 -30 3580 27
rect 3780 10 5510 27
rect 3780 -30 4220 10
rect 3568 -42 4220 -30
rect 3840 -200 4220 -42
rect 9770 -200 10210 830
rect 3840 -316 10210 -200
rect 1866 -484 10210 -316
rect 3840 -710 10210 -484
rect 3238 -1402 3248 -1321
rect 3472 -1402 3482 -1321
<< via1 >>
rect 3580 1667 3780 1724
rect 4000 1720 4081 1801
rect 5387 1717 5473 1803
rect 4640 1370 4700 1430
rect 4020 540 4080 600
rect 7560 1120 7650 1140
rect 7560 920 7577 1120
rect 7577 920 7634 1120
rect 7634 920 7650 1120
rect 7560 900 7650 920
rect 9400 860 10410 1120
rect 11464 905 11535 976
rect 4180 640 4240 700
rect 5270 640 5330 700
rect 5270 440 5330 500
rect 4640 130 4700 190
rect 3248 -1333 3472 -1321
rect 3248 -1390 3260 -1333
rect 3260 -1390 3460 -1333
rect 3460 -1390 3472 -1333
rect 3248 -1402 3472 -1390
<< metal2 >>
rect 3580 1724 3780 1734
rect 3994 1720 4000 1801
rect 4081 1720 4087 1801
rect 4643 1729 4703 1733
rect 4638 1724 4708 1729
rect 3580 1657 3780 1667
rect 4016 610 4065 1720
rect 4638 1664 4643 1724
rect 4703 1664 4708 1724
rect 5381 1717 5387 1803
rect 5473 1717 5479 1803
rect 4638 1430 4708 1664
rect 4638 1370 4640 1430
rect 4700 1370 4708 1430
rect 4638 1363 4708 1370
rect 4640 1360 4700 1363
rect 4180 700 4240 710
rect 5270 700 5330 710
rect 4240 650 5270 690
rect 4180 630 4240 640
rect 5270 630 5330 640
rect 4016 600 4080 610
rect 4016 540 4020 600
rect 4016 536 4080 540
rect 4020 530 4080 536
rect 5270 500 5330 510
rect 5408 493 5453 1717
rect 7560 1140 7650 1150
rect 7560 890 7650 900
rect 9400 1120 10410 1130
rect 11440 976 11560 1000
rect 11440 905 11464 976
rect 11535 905 11560 976
rect 11440 890 11560 905
rect 9400 850 10410 860
rect 5330 448 5453 493
rect 5270 430 5330 440
rect 4640 190 4700 200
rect 4634 130 4640 172
rect 4700 130 4716 172
rect 3248 -1320 3472 -1311
rect 4634 -1320 4716 130
rect 3248 -1321 4716 -1320
rect 3472 -1402 4716 -1321
rect 3248 -1412 3472 -1402
<< via2 >>
rect 3580 1667 3780 1724
rect 4643 1664 4703 1724
rect 7560 900 7650 1140
rect 9400 860 10410 1120
rect 11464 905 11535 976
<< metal3 >>
rect 3570 1724 4708 1729
rect 3570 1667 3580 1724
rect 3780 1667 4643 1724
rect 3570 1664 4643 1667
rect 4703 1664 4708 1724
rect 3570 1662 4708 1664
rect 3750 1659 4708 1662
rect 7550 1140 7660 1145
rect 7550 900 7560 1140
rect 7650 900 7660 1140
rect 7550 895 7660 900
rect 9390 1120 10420 1125
rect 9390 860 9400 1120
rect 10410 860 10420 1120
rect 11440 981 11560 1000
rect 11440 900 11459 981
rect 11540 900 11560 981
rect 11440 890 11560 900
rect 9390 855 10420 860
<< via3 >>
rect 7560 900 7650 1140
rect 9400 860 10410 1120
rect 11459 976 11540 981
rect 11459 905 11464 976
rect 11464 905 11535 976
rect 11535 905 11540 976
rect 11459 900 11540 905
<< metal4 >>
rect 7559 1140 7651 1141
rect 7559 900 7560 1140
rect 7650 900 7651 1140
rect 7559 899 7651 900
rect 9399 1120 10411 1121
rect 7560 640 7650 899
rect 9399 860 9400 1120
rect 10410 860 10411 1120
rect 11440 981 11560 1000
rect 11440 900 11459 981
rect 11540 900 11560 981
rect 11440 890 11560 900
rect 9399 859 10411 860
rect 9820 -1320 10100 859
rect 11464 525 11535 890
use sky130_fd_pr__res_generic_l1_3AQK6Q  R1
timestamp 1717183566
transform 0 1 6397 -1 0 1260
box -100 -877 100 877
use sky130_fd_pr__res_generic_l1_XY2C22  R2
timestamp 1717182944
transform 0 1 6577 -1 0 1020
box -100 -1057 100 1057
use sky130_fd_pr__res_generic_l1_3BGJFP  R4
timestamp 1717181420
transform 1 0 3360 0 1 307
box -100 -1697 100 1697
use sky130_fd_pr__nfet_01v8_BXYDM4  sky130_fd_pr__nfet_01v8_BXYDM4_0
timestamp 1717182944
transform 1 0 5301 0 1 289
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_NKKNMA  sky130_fd_pr__pfet_01v8_NKKNMA_0
timestamp 1717181835
transform 1 0 4881 0 1 1064
box -211 -484 211 484
use sky130_fd_pr__res_generic_l1_3AQK6Q  sky130_fd_pr__res_generic_l1_3AQK6Q_0
timestamp 1717183566
transform -1 0 3680 0 -1 847
box -100 -877 100 877
use sky130_fd_pr__cap_mim_m3_1_4PHTN9  XC1
timestamp 1717181420
transform -1 0 11196 0 1 -310
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_TNHPNJ  XC2
timestamp 1717182944
transform 1 0 7716 0 1 -310
box -2186 -1040 2186 1040
use sky130_fd_pr__pfet_01v8_GPKNM8  XM2
timestamp 1717182944
transform 1 0 5301 0 1 1064
box -211 -484 211 484
use sky130_fd_pr__nfet_01v8_BXYDM4  XM3
timestamp 1717182944
transform 1 0 4051 0 1 289
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_7P3MHC  XM4
timestamp 1717181835
transform 1 0 4051 0 1 964
box -211 -384 211 384
use sky130_fd_pr__nfet_01v8_5WP7M2  XM5
timestamp 1717181835
transform 1 0 4471 0 1 289
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_NKK3FE  XM8
timestamp 1717181835
transform 1 0 4461 0 1 1264
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_5WP7M2  XM9
timestamp 1717181835
transform 1 0 4881 0 1 289
box -211 -279 211 279
<< labels >>
flabel metal1 1850 1830 2050 2030 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 2250 1830 2450 2030 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 3940 1830 4140 2030 0 FreeSans 256 0 0 0 QA
port 2 nsew
flabel metal1 5330 1830 5530 2030 0 FreeSans 256 0 0 0 QB
port 3 nsew
flabel metal1 7990 1830 8190 2030 0 FreeSans 256 0 0 0 VOUT
port 4 nsew
<< end >>
