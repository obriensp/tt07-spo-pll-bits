magic
tech sky130A
magscale 1 2
timestamp 1717026976
<< pwell >>
rect -241 -279 241 279
<< nmos >>
rect -45 -131 45 69
<< ndiff >>
rect -103 57 -45 69
rect -103 -119 -91 57
rect -57 -119 -45 57
rect -103 -131 -45 -119
rect 45 57 103 69
rect 45 -119 57 57
rect 91 -119 103 57
rect 45 -131 103 -119
<< ndiffc >>
rect -91 -119 -57 57
rect 57 -119 91 57
<< psubdiff >>
rect -205 209 -109 243
rect 109 209 205 243
rect -205 147 -171 209
rect 171 147 205 209
rect -205 -209 -171 -147
rect 171 -209 205 -147
rect -205 -243 -109 -209
rect 109 -243 205 -209
<< psubdiffcont >>
rect -109 209 109 243
rect -205 -147 -171 147
rect 171 -147 205 147
rect -109 -243 109 -209
<< poly >>
rect -45 141 45 157
rect -45 107 -29 141
rect 29 107 45 141
rect -45 69 45 107
rect -45 -157 45 -131
<< polycont >>
rect -29 107 29 141
<< locali >>
rect -125 209 -109 243
rect 109 209 125 243
rect -205 147 -171 163
rect 171 147 205 163
rect -45 107 -29 141
rect 29 107 45 141
rect -91 57 -57 73
rect -91 -135 -57 -119
rect 57 57 91 73
rect 57 -135 91 -119
rect -205 -163 -171 -147
rect 171 -163 205 -147
rect -125 -243 -109 -209
rect 109 -243 125 -209
<< viali >>
rect -29 107 29 141
rect -91 -119 -57 57
rect 57 -119 91 57
<< metal1 >>
rect -41 141 41 147
rect -41 107 -29 141
rect 29 107 41 141
rect -41 101 41 107
rect -97 57 -51 69
rect -97 -119 -91 57
rect -57 -119 -51 57
rect -97 -131 -51 -119
rect 51 57 97 69
rect 51 -119 57 57
rect 91 -119 97 57
rect 51 -131 97 -119
<< properties >>
string FIXED_BBOX -188 -226 188 226
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.45 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
