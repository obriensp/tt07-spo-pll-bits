magic
tech sky130A
magscale 1 2
timestamp 1717119155
<< viali >>
rect 2136 1731 2170 1969
rect 2771 1862 2805 1896
rect 2949 1862 2983 1896
rect 3046 1862 3080 1896
rect 3332 1794 3366 1828
rect 3792 1799 3826 1901
rect 3976 1799 4010 1901
rect -94 1154 4 1252
rect -68 393 -34 895
rect -68 -888 -34 -394
rect -514 -1194 -416 -1096
<< metal1 >>
rect -530 2080 -520 2170
rect -410 2080 2170 2170
rect 2124 1969 2182 1981
rect 710 1800 720 1870
rect 780 1849 790 1870
rect 2124 1849 2136 1969
rect 780 1820 2136 1849
rect 780 1800 790 1820
rect 2124 1731 2136 1820
rect 2170 1731 2182 1969
rect 2753 1850 2763 1908
rect 2821 1850 2831 1908
rect 2908 1850 2918 1910
rect 2976 1896 2995 1910
rect 2983 1862 2995 1896
rect 2976 1850 2995 1862
rect 3024 1850 3034 1910
rect 3092 1850 3102 1910
rect 3780 1902 3838 1913
rect 3768 1901 3850 1902
rect 3768 1896 3792 1901
rect 3826 1896 3850 1901
rect 3320 1839 3378 1842
rect 3320 1787 3330 1839
rect 3382 1787 3388 1839
rect 3768 1826 3774 1896
rect 3844 1826 3850 1896
rect 3964 1901 4022 1913
rect 3964 1881 3976 1901
rect 3768 1820 3792 1826
rect 3780 1799 3792 1820
rect 3826 1820 3850 1826
rect 3949 1875 3976 1881
rect 4010 1881 4022 1901
rect 4010 1875 4031 1881
rect 3826 1799 3838 1820
rect 3949 1805 3955 1875
rect 4025 1805 4031 1875
rect 3949 1799 3976 1805
rect 4010 1799 4031 1805
rect 3780 1787 3838 1799
rect 3964 1787 4022 1799
rect 3320 1783 3378 1787
rect 2124 1719 2182 1731
rect -110 1530 -100 1620
rect 10 1530 2170 1620
rect -106 1260 16 1264
rect -460 1258 4590 1260
rect -460 1150 -100 1258
rect -110 1148 -100 1150
rect 10 1150 4590 1258
rect 10 1148 16 1150
rect -110 1142 16 1148
rect -110 895 -20 1142
rect -110 880 -68 895
rect -310 440 -250 880
rect -190 480 -68 880
rect -310 350 -190 440
rect -110 393 -68 480
rect -34 393 -20 895
rect 160 580 170 650
rect 330 580 340 650
rect 670 580 680 650
rect 840 580 850 650
rect 1180 580 1190 650
rect 1350 580 1360 650
rect 1690 580 1700 650
rect 1860 580 1870 650
rect 2200 580 2210 650
rect 2370 580 2380 650
rect 2710 580 2720 650
rect 2880 580 2890 650
rect 3220 580 3230 650
rect 3390 580 3400 650
rect -110 380 -20 393
rect -310 180 -250 350
rect -340 80 -330 180
rect -230 80 -220 180
rect -310 -800 -250 80
rect 30 -240 40 -130
rect 190 -240 200 -130
rect 1370 -240 1380 -130
rect 1530 -240 1540 -130
rect 2390 -240 2400 -130
rect 2550 -240 2560 -130
rect 3410 -240 3420 -130
rect 3570 -240 3580 -130
rect 4430 -240 4440 -130
rect 4590 -240 4600 -130
rect -90 -394 -20 -380
rect -90 -420 -68 -394
rect -190 -800 -68 -420
rect -280 -930 -270 -840
rect -180 -930 -170 -840
rect -90 -888 -68 -800
rect -34 -888 -20 -394
rect 160 -800 170 -730
rect 330 -800 340 -730
rect 670 -800 680 -730
rect 840 -800 850 -730
rect 1180 -800 1190 -730
rect 1350 -800 1360 -730
rect 1690 -800 1700 -730
rect 1860 -800 1870 -730
rect 2200 -800 2210 -730
rect 2370 -800 2380 -730
rect 2710 -800 2720 -730
rect 2880 -800 2890 -730
rect 3220 -800 3230 -730
rect 3390 -800 3400 -730
rect -526 -1090 -404 -1084
rect -90 -1090 -20 -888
rect -526 -1200 -520 -1090
rect -410 -1200 4590 -1090
rect -526 -1206 -404 -1200
<< via1 >>
rect -520 2080 -410 2170
rect 720 1800 780 1870
rect 2763 1896 2821 1908
rect 2763 1862 2771 1896
rect 2771 1862 2805 1896
rect 2805 1862 2821 1896
rect 2763 1850 2821 1862
rect 2918 1896 2976 1910
rect 2918 1862 2949 1896
rect 2949 1862 2976 1896
rect 2918 1850 2976 1862
rect 3034 1896 3092 1910
rect 3034 1862 3046 1896
rect 3046 1862 3080 1896
rect 3080 1862 3092 1896
rect 3034 1850 3092 1862
rect 3330 1828 3382 1839
rect 3330 1794 3332 1828
rect 3332 1794 3366 1828
rect 3366 1794 3382 1828
rect 3330 1787 3382 1794
rect 3774 1826 3792 1896
rect 3792 1826 3826 1896
rect 3826 1826 3844 1896
rect 3955 1805 3976 1875
rect 3976 1805 4010 1875
rect 4010 1805 4025 1875
rect -100 1530 10 1620
rect -100 1252 10 1258
rect -100 1154 -94 1252
rect -94 1154 4 1252
rect 4 1154 10 1252
rect -100 1148 10 1154
rect 170 580 330 650
rect 680 580 840 650
rect 1190 580 1350 650
rect 1700 580 1860 650
rect 2210 580 2370 650
rect 2720 580 2880 650
rect 3230 580 3390 650
rect 3740 580 3900 650
rect 4250 580 4410 650
rect -330 80 -230 180
rect 40 -240 190 -130
rect 1380 -240 1530 -130
rect 2400 -240 2550 -130
rect 3420 -240 3570 -130
rect 4440 -240 4590 -130
rect -270 -930 -180 -840
rect 170 -800 330 -730
rect 680 -800 840 -730
rect 1190 -800 1350 -730
rect 1700 -800 1860 -730
rect 2210 -800 2370 -730
rect 2720 -800 2880 -730
rect 3230 -800 3390 -730
rect 3740 -800 3900 -730
rect 4250 -800 4410 -730
rect -520 -1096 -410 -1090
rect -520 -1194 -514 -1096
rect -514 -1194 -416 -1096
rect -416 -1194 -410 -1096
rect -520 -1200 -410 -1194
<< metal2 >>
rect 1096 2190 1214 2199
rect -520 2170 -410 2180
rect 1096 2090 1105 2190
rect 1205 2090 1214 2190
rect 1096 2081 1214 2090
rect -520 2070 -410 2080
rect 720 1870 780 1880
rect 720 1790 780 1800
rect -100 1620 10 1630
rect -100 1520 10 1530
rect 1131 1301 1180 2081
rect 1496 2062 1505 2162
rect 1605 2062 1614 2162
rect 1530 1907 1581 2062
rect 2763 1908 2821 1918
rect 1530 1856 2763 1907
rect 2763 1840 2821 1850
rect 2918 1910 2976 1920
rect 2918 1840 2976 1850
rect 3034 1910 3092 1920
rect 3034 1840 3092 1850
rect 3768 1896 3850 1902
rect 2921 1403 2970 1840
rect 3039 1556 3086 1840
rect 3330 1839 3382 1845
rect 3768 1826 3774 1896
rect 3844 1826 3850 1896
rect 3768 1820 3850 1826
rect 3949 1875 4031 1881
rect 3949 1805 3955 1875
rect 4025 1805 4031 1875
rect 3949 1799 4031 1805
rect 3330 1781 3382 1787
rect 3032 1547 3092 1556
rect 3032 1478 3092 1487
rect 2906 1343 2915 1403
rect 2975 1343 2984 1403
rect 3331 1301 3380 1781
rect -106 1258 16 1264
rect -106 1148 -100 1258
rect 10 1148 16 1258
rect 1131 1252 3380 1301
rect -106 1142 16 1148
rect -330 650 4590 670
rect -330 580 170 650
rect 330 580 680 650
rect 840 580 1190 650
rect 1350 580 1700 650
rect 1860 580 2210 650
rect 2370 580 2720 650
rect 2880 580 3230 650
rect 3390 580 3740 650
rect 3900 580 4250 650
rect 4410 580 4590 650
rect -330 560 4590 580
rect -330 180 -230 560
rect -129 219 -29 223
rect -330 70 -230 80
rect -134 214 -24 219
rect -134 114 -129 214
rect -29 114 -24 214
rect -134 -730 -24 114
rect 40 -130 190 -120
rect 40 -250 190 -240
rect 1380 -130 1530 -120
rect 1380 -250 1530 -240
rect 2400 -130 2550 -120
rect 2400 -250 2550 -240
rect 3420 -130 3570 -120
rect 3420 -250 3570 -240
rect 4440 -130 4590 -120
rect 4440 -250 4590 -240
rect 150 -730 4590 -710
rect -460 -800 170 -730
rect 330 -800 680 -730
rect 840 -800 1190 -730
rect 1350 -800 1700 -730
rect 1860 -800 2210 -730
rect 2370 -800 2720 -730
rect 2880 -800 3230 -730
rect 3390 -800 3740 -730
rect 3900 -800 4250 -730
rect 4410 -800 4590 -730
rect -270 -840 -180 -800
rect 150 -820 4590 -800
rect -270 -940 -180 -930
rect -526 -1090 -404 -1084
rect -526 -1200 -520 -1090
rect -410 -1200 -404 -1090
rect -526 -1206 -404 -1200
<< via2 >>
rect -520 2080 -410 2170
rect 1105 2090 1205 2190
rect 720 1800 780 1870
rect -100 1530 10 1620
rect 1505 2062 1605 2162
rect 3779 1831 3839 1891
rect 3960 1810 4020 1870
rect 3032 1487 3092 1547
rect 2915 1343 2975 1403
rect -95 1153 5 1253
rect -129 114 -29 214
rect 40 -240 190 -130
rect 1380 -240 1530 -130
rect 2400 -240 2550 -130
rect 3420 -240 3570 -130
rect 4440 -240 4590 -130
rect -515 -1195 -415 -1095
<< metal3 >>
rect -520 2175 -410 2230
rect -530 2170 -400 2175
rect -530 2080 -520 2170
rect -410 2080 -400 2170
rect -530 2075 -400 2080
rect -520 -1095 -410 2075
rect -100 1625 10 2230
rect -110 1620 20 1625
rect -110 1530 -100 1620
rect 10 1530 20 1620
rect -110 1525 20 1530
rect -100 1253 10 1525
rect -100 1153 -95 1253
rect 5 1153 10 1253
rect -100 1148 10 1153
rect 310 219 420 2230
rect 700 2030 810 2230
rect 1100 2190 1210 2230
rect 1100 2090 1105 2190
rect 1205 2090 1210 2190
rect 1100 2030 1210 2090
rect 1500 2162 1610 2230
rect 1500 2062 1505 2162
rect 1605 2062 1610 2162
rect 1500 2030 1610 2062
rect 3470 2035 4025 2105
rect 719 1875 784 2030
rect 710 1870 790 1875
rect 710 1800 720 1870
rect 780 1800 790 1870
rect 710 1795 790 1800
rect -134 214 420 219
rect -134 114 -129 214
rect -29 114 420 214
rect -134 109 420 114
rect 30 -130 200 -125
rect 30 -240 40 -130
rect 190 -146 200 -130
rect 719 -146 784 1795
rect 1420 1547 3097 1552
rect 1420 1487 3032 1547
rect 3092 1487 3097 1547
rect 1420 1482 3097 1487
rect 1420 -125 1490 1482
rect 2440 1403 2980 1408
rect 2440 1343 2915 1403
rect 2975 1343 2980 1403
rect 2440 1338 2980 1343
rect 2440 -125 2510 1338
rect 3470 -125 3540 2035
rect 3774 1891 3844 1896
rect 3774 1831 3779 1891
rect 3839 1831 3844 1891
rect 3774 1434 3844 1831
rect 3955 1870 4025 2035
rect 3955 1810 3960 1870
rect 4020 1810 4025 1870
rect 3955 1805 4025 1810
rect 3774 1364 4560 1434
rect 4490 -125 4560 1364
rect 190 -211 784 -146
rect 1370 -130 1540 -125
rect 190 -240 200 -211
rect 30 -245 200 -240
rect 1370 -240 1380 -130
rect 1530 -240 1540 -130
rect 1370 -245 1540 -240
rect 2390 -130 2560 -125
rect 2390 -240 2400 -130
rect 2550 -240 2560 -130
rect 2390 -245 2560 -240
rect 3410 -130 3580 -125
rect 3410 -240 3420 -130
rect 3570 -240 3580 -130
rect 3410 -245 3580 -240
rect 4430 -130 4600 -125
rect 4430 -240 4440 -130
rect 4590 -240 4600 -130
rect 4430 -245 4600 -240
rect -520 -1195 -515 -1095
rect -415 -1195 -410 -1095
rect -520 -1200 -410 -1195
use delay_stage  delay_stage_0 ~/Development/spo/vlsi/tt07-spo-pll/mag
timestamp 1717029282
transform 1 0 -90 0 1 1470
box 1110 -2670 1620 -210
use delay_stage  delay_stage_1
timestamp 1717029282
transform 1 0 2970 0 1 1470
box 1110 -2670 1620 -210
use delay_stage  delay_stage_2
timestamp 1717029282
transform 1 0 1440 0 1 1470
box 1110 -2670 1620 -210
use delay_stage  delay_stage_3
timestamp 1717029282
transform 1 0 2460 0 1 1470
box 1110 -2670 1620 -210
use delay_stage  delay_stage_4
timestamp 1717029282
transform 1 0 930 0 1 1470
box 1110 -2670 1620 -210
use delay_stage  delay_stage_5
timestamp 1717029282
transform 1 0 420 0 1 1470
box 1110 -2670 1620 -210
use delay_stage  delay_stage_6
timestamp 1717029282
transform 1 0 1950 0 1 1470
box 1110 -2670 1620 -210
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_0
timestamp 1704896540
transform -1 0 4040 0 -1 2122
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1704896540
transform -1 0 4132 0 -1 2122
box -38 -48 130 592
use delay_stage  x1
timestamp 1717029282
transform 1 0 -1110 0 1 1470
box 1110 -2670 1620 -210
use delay_stage  x2
timestamp 1717029282
transform 1 0 -600 0 1 1470
box 1110 -2670 1620 -210
use sky130_fd_pr__pfet_01v8_PLD8WZ  XM5
timestamp 1717055118
transform 1 0 -224 0 1 644
box -226 -384 226 384
use sky130_fd_pr__nfet_01v8_lvt_TKZJHP  XM6
timestamp 1717055118
transform 1 0 -224 0 1 -641
box -226 -379 226 379
<< labels >>
flabel metal3 -520 2030 -410 2230 0 FreeSans 160 0 0 0 vss
port 0 nsew
flabel metal3 -100 2030 10 2230 0 FreeSans 160 0 0 0 vdd
port 1 nsew
flabel metal3 310 2030 420 2230 0 FreeSans 160 0 0 0 vcont
port 2 nsew
flabel metal3 700 2030 810 2230 0 FreeSans 160 0 0 0 out
port 3 nsew
flabel metal3 1100 2030 1210 2230 0 FreeSans 160 0 0 0 s0
port 4 nsew
flabel metal3 1500 2030 1610 2230 0 FreeSans 160 0 0 0 s1
port 5 nsew
<< end >>
