magic
tech sky130A
magscale 1 2
timestamp 1717208985
<< viali >>
rect 1232 -222 1390 -188
rect 1652 -222 1810 -188
rect 2072 -222 2230 -188
rect 2492 -222 2650 -188
rect 1232 -1464 1390 -1430
rect 1652 -1464 1810 -1430
rect 2072 -1464 2230 -1430
rect 2492 -1464 2650 -1430
<< metal1 >>
rect 800 -160 2800 -140
rect 800 -188 1470 -160
rect 800 -222 1232 -188
rect 1390 -220 1470 -188
rect 1530 -188 2800 -160
rect 1530 -220 1652 -188
rect 1390 -222 1652 -220
rect 1810 -222 2072 -188
rect 2230 -222 2492 -188
rect 2650 -222 2800 -188
rect 800 -240 2800 -222
rect 800 -340 1000 -240
rect 1034 -340 1040 -280
rect 1100 -340 1350 -280
rect 800 -877 1000 -810
rect 800 -963 847 -877
rect 933 -880 1000 -877
rect 1240 -880 1290 -380
rect 933 -950 1290 -880
rect 933 -963 1000 -950
rect 800 -1010 1000 -963
rect 1240 -1280 1290 -950
rect 1330 -900 1380 -380
rect 1630 -700 1710 -240
rect 1750 -700 1910 -300
rect 2050 -700 2130 -240
rect 2170 -700 2330 -300
rect 2470 -700 2550 -240
rect 2590 -500 2750 -300
rect 2800 -500 3000 -450
rect 2590 -610 3000 -500
rect 2590 -700 2750 -610
rect 2800 -650 3000 -610
rect 1700 -900 1760 -740
rect 1330 -950 1760 -900
rect 1330 -1280 1380 -950
rect 1700 -1120 1760 -950
rect 1860 -1050 1910 -700
rect 2120 -880 2180 -740
rect 2090 -970 2100 -880
rect 2190 -970 2200 -880
rect 2280 -890 2330 -700
rect 2540 -890 2600 -740
rect 2280 -950 2600 -890
rect 1840 -1130 1850 -1050
rect 1930 -1130 1940 -1050
rect 2120 -1120 2180 -970
rect 1840 -1150 1910 -1130
rect 2280 -1150 2330 -950
rect 2540 -1120 2600 -950
rect 2700 -1150 2750 -700
rect 1470 -1320 1530 -1314
rect 800 -1420 1000 -1320
rect 1280 -1380 1470 -1320
rect 1470 -1386 1530 -1380
rect 1630 -1420 1710 -1150
rect 1750 -1360 1910 -1150
rect 2050 -1420 2130 -1150
rect 2170 -1360 2330 -1150
rect 2470 -1420 2550 -1150
rect 2590 -1360 2750 -1150
rect 2800 -1048 3000 -990
rect 2800 -1142 2863 -1048
rect 2957 -1142 3000 -1048
rect 2800 -1190 3000 -1142
rect 800 -1430 2800 -1420
rect 800 -1490 1040 -1430
rect 1100 -1464 1232 -1430
rect 1390 -1464 1652 -1430
rect 1810 -1464 2072 -1430
rect 2230 -1464 2492 -1430
rect 2650 -1464 2800 -1430
rect 1100 -1490 2800 -1464
rect 800 -1520 2800 -1490
<< via1 >>
rect 1470 -220 1530 -160
rect 1040 -340 1100 -280
rect 847 -963 933 -877
rect 2100 -970 2190 -880
rect 1850 -1130 1930 -1050
rect 1470 -1380 1530 -1320
rect 2863 -1142 2957 -1048
rect 1040 -1490 1100 -1430
<< metal2 >>
rect 1460 -160 1540 -150
rect 1460 -220 1470 -160
rect 1530 -220 1540 -160
rect 1460 -230 1540 -220
rect 1030 -280 1110 -270
rect 1030 -340 1040 -280
rect 1100 -340 1110 -280
rect 1030 -350 1110 -340
rect 847 -877 933 -871
rect 2100 -880 2190 -870
rect 933 -948 2100 -892
rect 2070 -950 2100 -948
rect 847 -969 933 -963
rect 2100 -980 2190 -970
rect 1850 -1050 1930 -1040
rect 2850 -1048 2970 -1040
rect 2850 -1070 2863 -1048
rect 1930 -1120 2863 -1070
rect 1850 -1140 1930 -1130
rect 2850 -1142 2863 -1120
rect 2957 -1142 2970 -1048
rect 2850 -1150 2970 -1142
rect 1460 -1320 1540 -1310
rect 1460 -1380 1470 -1320
rect 1530 -1380 1540 -1320
rect 1460 -1390 1540 -1380
rect 1030 -1430 1110 -1420
rect 1030 -1490 1040 -1430
rect 1100 -1490 1110 -1430
rect 1030 -1500 1110 -1490
<< via2 >>
rect 1472 -218 1528 -162
rect 1040 -340 1100 -280
rect 1470 -1380 1530 -1320
rect 1042 -1488 1098 -1432
<< metal3 >>
rect 1467 -162 1533 -157
rect 1467 -218 1472 -162
rect 1528 -218 1533 -162
rect 1467 -223 1533 -218
rect 1035 -280 1105 -275
rect 1035 -340 1040 -280
rect 1100 -340 1105 -280
rect 1035 -345 1105 -340
rect 1040 -1427 1100 -345
rect 1470 -1315 1530 -223
rect 1465 -1320 1535 -1315
rect 1465 -1380 1470 -1320
rect 1530 -1380 1535 -1320
rect 1465 -1385 1535 -1380
rect 1037 -1432 1103 -1427
rect 1037 -1488 1042 -1432
rect 1098 -1488 1103 -1432
rect 1037 -1493 1103 -1488
use sky130_fd_pr__nfet_01v8_BXYDM4  sky130_fd_pr__nfet_01v8_BXYDM4_0
timestamp 1717207579
transform 1 0 2571 0 1 -1221
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_7P3MHC  sky130_fd_pr__pfet_01v8_7P3MHC_0
timestamp 1717207579
transform 1 0 2571 0 1 -536
box -211 -384 211 384
use sky130_fd_pr__nfet_01v8_BXYDM4  XM1
timestamp 1717207579
transform 1 0 2151 0 1 -1221
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_7P3MHC  XM4
timestamp 1717207579
transform 1 0 2151 0 1 -536
box -211 -384 211 384
use sky130_fd_pr__nfet_01v8_5WP7M2  XM5
timestamp 1717207579
transform 1 0 1311 0 1 -1221
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_NK3MHE  XM6
timestamp 1717207579
transform 1 0 1311 0 1 -536
box -211 -384 211 384
use sky130_fd_pr__nfet_01v8_BXYDM4  XM7
timestamp 1717207579
transform 1 0 1731 0 1 -1221
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_7P3MHC  XM8
timestamp 1717207579
transform 1 0 1731 0 1 -536
box -211 -384 211 384
<< labels >>
flabel metal1 800 -1520 1000 -1320 0 FreeSans 256 0 0 0 vss
port 4 nsew
flabel metal1 800 -340 1000 -140 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 2800 -1190 3000 -990 0 FreeSans 256 0 0 0 clk_inverted
port 3 nsew
flabel metal1 2800 -650 3000 -450 0 FreeSans 256 0 0 0 clk_delayed
port 1 nsew
flabel metal1 800 -1010 1000 -810 0 FreeSans 256 0 0 0 clk
port 2 nsew
<< end >>
