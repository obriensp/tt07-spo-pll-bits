magic
tech sky130A
magscale 1 2
timestamp 1717181420
<< locali >>
rect -100 1640 100 1697
rect -100 -1697 100 -1640
<< rlocali >>
rect -100 -1640 100 1640
<< properties >>
string gencell sky130_fd_pr__res_generic_l1
string library sky130
string parameters w 1.0 l 16.4 m 1 nx 1 wmin 0.17 lmin 0.17 rho 12.8 val 209.92 dummy 0 dw 0.0 term 0.0 snake 0 roverlap 0
<< end >>
