magic
tech sky130A
magscale 1 2
timestamp 1716920833
<< viali >>
rect 2237 9537 2271 9571
rect 2421 9469 2455 9503
rect 3249 9469 3283 9503
rect 3709 9469 3743 9503
rect 5181 9469 5215 9503
rect 5641 9469 5675 9503
rect 6009 9469 6043 9503
rect 6101 9469 6135 9503
rect 6377 9469 6411 9503
rect 7297 9469 7331 9503
rect 7481 9469 7515 9503
rect 8401 9469 8435 9503
rect 1970 9401 2004 9435
rect 4936 9401 4970 9435
rect 8646 9401 8680 9435
rect 857 9333 891 9367
rect 3065 9333 3099 9367
rect 3433 9333 3467 9367
rect 3525 9333 3559 9367
rect 3801 9333 3835 9367
rect 5457 9333 5491 9367
rect 5825 9333 5859 9367
rect 6285 9333 6319 9367
rect 7021 9333 7055 9367
rect 7113 9333 7147 9367
rect 8125 9333 8159 9367
rect 9781 9333 9815 9367
rect 1593 9129 1627 9163
rect 5641 9129 5675 9163
rect 7205 9129 7239 9163
rect 9689 9129 9723 9163
rect 2728 9061 2762 9095
rect 4528 9061 4562 9095
rect 7564 9061 7598 9095
rect 857 8993 891 9027
rect 3249 8993 3283 9027
rect 4261 8993 4295 9027
rect 5825 8993 5859 9027
rect 6092 8993 6126 9027
rect 7297 8993 7331 9027
rect 9505 8993 9539 9027
rect 2973 8925 3007 8959
rect 3617 8925 3651 8959
rect 9413 8925 9447 8959
rect 8769 8857 8803 8891
rect 1501 8789 1535 8823
rect 3065 8789 3099 8823
rect 4169 8789 4203 8823
rect 8677 8789 8711 8823
rect 1501 8585 1535 8619
rect 4629 8585 4663 8619
rect 6745 8585 6779 8619
rect 9781 8585 9815 8619
rect 6193 8517 6227 8551
rect 4813 8449 4847 8483
rect 6837 8449 6871 8483
rect 857 8381 891 8415
rect 1317 8381 1351 8415
rect 1593 8381 1627 8415
rect 3249 8381 3283 8415
rect 5069 8381 5103 8415
rect 6561 8381 6595 8415
rect 8401 8381 8435 8415
rect 1838 8313 1872 8347
rect 3494 8313 3528 8347
rect 7104 8313 7138 8347
rect 8646 8313 8680 8347
rect 1041 8245 1075 8279
rect 2973 8245 3007 8279
rect 8217 8245 8251 8279
rect 2697 8041 2731 8075
rect 8677 8041 8711 8075
rect 3985 7905 4019 7939
rect 6949 7905 6983 7939
rect 7205 7905 7239 7939
rect 7389 7905 7423 7939
rect 9781 7905 9815 7939
rect 5825 7701 5859 7735
rect 9229 7701 9263 7735
rect 8125 7497 8159 7531
rect 4629 7429 4663 7463
rect 3249 7361 3283 7395
rect 5273 7361 5307 7395
rect 7849 7361 7883 7395
rect 857 7293 891 7327
rect 1124 7293 1158 7327
rect 3505 7293 3539 7327
rect 6009 7293 6043 7327
rect 7593 7293 7627 7327
rect 7941 7293 7975 7327
rect 9873 7293 9907 7327
rect 9606 7225 9640 7259
rect 2237 7157 2271 7191
rect 4721 7157 4755 7191
rect 6101 7157 6135 7191
rect 6469 7157 6503 7191
rect 8493 7157 8527 7191
rect 8524 6885 8558 6919
rect 1981 6817 2015 6851
rect 2881 6817 2915 6851
rect 3884 6817 3918 6851
rect 8769 6817 8803 6851
rect 9505 6817 9539 6851
rect 9873 6817 9907 6851
rect 2237 6749 2271 6783
rect 3617 6749 3651 6783
rect 9689 6681 9723 6715
rect 857 6613 891 6647
rect 2329 6613 2363 6647
rect 4997 6613 5031 6647
rect 7389 6613 7423 6647
rect 8861 6613 8895 6647
rect 3801 6409 3835 6443
rect 9781 6409 9815 6443
rect 4353 6341 4387 6375
rect 7113 6341 7147 6375
rect 7757 6341 7791 6375
rect 949 6273 983 6307
rect 3525 6273 3559 6307
rect 5733 6273 5767 6307
rect 8401 6273 8435 6307
rect 1685 6205 1719 6239
rect 3433 6205 3467 6239
rect 6101 6205 6135 6239
rect 6377 6205 6411 6239
rect 6561 6205 6595 6239
rect 6837 6205 6871 6239
rect 7297 6205 7331 6239
rect 7389 6205 7423 6239
rect 7481 6205 7515 6239
rect 8657 6205 8691 6239
rect 1593 6137 1627 6171
rect 1930 6137 1964 6171
rect 5488 6137 5522 6171
rect 5825 6137 5859 6171
rect 6653 6137 6687 6171
rect 7113 6137 7147 6171
rect 7757 6137 7791 6171
rect 3065 6069 3099 6103
rect 5923 6069 5957 6103
rect 6009 6069 6043 6103
rect 6561 6069 6595 6103
rect 7021 6069 7055 6103
rect 7573 6069 7607 6103
rect 5549 5865 5583 5899
rect 6738 5865 6772 5899
rect 9137 5865 9171 5899
rect 9229 5865 9263 5899
rect 2136 5797 2170 5831
rect 6469 5797 6503 5831
rect 7297 5797 7331 5831
rect 4445 5729 4479 5763
rect 4905 5729 4939 5763
rect 6285 5729 6319 5763
rect 6561 5729 6595 5763
rect 6653 5729 6687 5763
rect 6837 5729 6871 5763
rect 7205 5729 7239 5763
rect 7757 5729 7791 5763
rect 8013 5729 8047 5763
rect 9781 5729 9815 5763
rect 1869 5661 1903 5695
rect 4261 5661 4295 5695
rect 4813 5661 4847 5695
rect 5825 5661 5859 5695
rect 6193 5661 6227 5695
rect 7021 5661 7055 5695
rect 4721 5593 4755 5627
rect 7665 5593 7699 5627
rect 3249 5525 3283 5559
rect 8401 5321 8435 5355
rect 6561 5185 6595 5219
rect 9045 5185 9079 5219
rect 3249 5117 3283 5151
rect 3433 5117 3467 5151
rect 6653 5117 6687 5151
rect 6837 5117 6871 5151
rect 2697 5049 2731 5083
rect 2881 5049 2915 5083
rect 3341 5049 3375 5083
rect 4813 5049 4847 5083
rect 7021 5049 7055 5083
rect 2513 4981 2547 5015
rect 4169 4777 4203 4811
rect 4905 4777 4939 4811
rect 5457 4777 5491 4811
rect 6929 4777 6963 4811
rect 7021 4777 7055 4811
rect 7389 4777 7423 4811
rect 2697 4709 2731 4743
rect 3801 4709 3835 4743
rect 3985 4709 4019 4743
rect 4537 4709 4571 4743
rect 4629 4709 4663 4743
rect 6837 4709 6871 4743
rect 949 4641 983 4675
rect 1216 4641 1250 4675
rect 2513 4641 2547 4675
rect 3249 4641 3283 4675
rect 4261 4641 4295 4675
rect 4409 4641 4443 4675
rect 4765 4641 4799 4675
rect 5516 4641 5550 4675
rect 5825 4641 5859 4675
rect 6009 4641 6043 4675
rect 6101 4641 6135 4675
rect 6377 4641 6411 4675
rect 7757 4641 7791 4675
rect 9137 4641 9171 4675
rect 3341 4573 3375 4607
rect 3617 4573 3651 4607
rect 4997 4573 5031 4607
rect 6193 4573 6227 4607
rect 7849 4573 7883 4607
rect 9229 4573 9263 4607
rect 2329 4505 2363 4539
rect 5641 4505 5675 4539
rect 6561 4505 6595 4539
rect 7205 4505 7239 4539
rect 8769 4505 8803 4539
rect 2881 4437 2915 4471
rect 5089 4437 5123 4471
rect 6653 4437 6687 4471
rect 2881 4233 2915 4267
rect 8861 4233 8895 4267
rect 7665 4165 7699 4199
rect 3341 4097 3375 4131
rect 7849 4097 7883 4131
rect 9045 4097 9079 4131
rect 1225 4029 1259 4063
rect 3249 4029 3283 4063
rect 3433 4029 3467 4063
rect 5273 4029 5307 4063
rect 5641 4029 5675 4063
rect 5825 4029 5859 4063
rect 6009 4029 6043 4063
rect 6101 4029 6135 4063
rect 6193 4029 6227 4063
rect 6377 4029 6411 4063
rect 6469 4029 6503 4063
rect 7021 4029 7055 4063
rect 7205 4029 7239 4063
rect 7297 4029 7331 4063
rect 7481 4029 7515 4063
rect 7757 4029 7791 4063
rect 9137 4029 9171 4063
rect 1492 3961 1526 3995
rect 2865 3961 2899 3995
rect 3065 3961 3099 3995
rect 2605 3893 2639 3927
rect 2697 3893 2731 3927
rect 3985 3893 4019 3927
rect 2053 3689 2087 3723
rect 2303 3689 2337 3723
rect 3157 3689 3191 3723
rect 3433 3689 3467 3723
rect 3801 3689 3835 3723
rect 5917 3689 5951 3723
rect 8953 3689 8987 3723
rect 2513 3621 2547 3655
rect 3525 3621 3559 3655
rect 3985 3621 4019 3655
rect 4528 3621 4562 3655
rect 7665 3621 7699 3655
rect 1869 3553 1903 3587
rect 2053 3553 2087 3587
rect 2973 3553 3007 3587
rect 3617 3553 3651 3587
rect 3893 3553 3927 3587
rect 6009 3553 6043 3587
rect 6929 3553 6963 3587
rect 7113 3553 7147 3587
rect 7205 3553 7239 3587
rect 7297 3553 7331 3587
rect 2697 3485 2731 3519
rect 2789 3485 2823 3519
rect 2881 3485 2915 3519
rect 4261 3485 4295 3519
rect 2145 3417 2179 3451
rect 3249 3417 3283 3451
rect 5641 3417 5675 3451
rect 2329 3349 2363 3383
rect 7573 3349 7607 3383
rect 4629 3145 4663 3179
rect 5457 3145 5491 3179
rect 7665 3145 7699 3179
rect 8033 3145 8067 3179
rect 9781 3145 9815 3179
rect 4813 3077 4847 3111
rect 8401 3009 8435 3043
rect 3249 2941 3283 2975
rect 4721 2941 4755 2975
rect 7573 2941 7607 2975
rect 7757 2941 7791 2975
rect 8657 2941 8691 2975
rect 3516 2873 3550 2907
rect 5273 2873 5307 2907
rect 5473 2873 5507 2907
rect 8217 2873 8251 2907
rect 5641 2805 5675 2839
rect 7849 2805 7883 2839
rect 8017 2805 8051 2839
rect 3525 2601 3559 2635
rect 5273 2601 5307 2635
rect 6193 2601 6227 2635
rect 7481 2601 7515 2635
rect 9505 2601 9539 2635
rect 3677 2533 3711 2567
rect 3893 2533 3927 2567
rect 5917 2533 5951 2567
rect 7113 2533 7147 2567
rect 7329 2533 7363 2567
rect 7941 2533 7975 2567
rect 8392 2533 8426 2567
rect 5089 2465 5123 2499
rect 5365 2465 5399 2499
rect 5641 2465 5675 2499
rect 6101 2465 6135 2499
rect 6285 2465 6319 2499
rect 6469 2465 6503 2499
rect 7021 2465 7055 2499
rect 7757 2465 7791 2499
rect 8033 2465 8067 2499
rect 8125 2465 8159 2499
rect 7573 2329 7607 2363
rect 3709 2261 3743 2295
rect 4905 2261 4939 2295
rect 5549 2261 5583 2295
rect 6929 2261 6963 2295
rect 7297 2261 7331 2295
rect 5641 2057 5675 2091
rect 6285 2057 6319 2091
rect 6561 2057 6595 2091
rect 8493 2057 8527 2091
rect 8769 2057 8803 2091
rect 4261 1921 4295 1955
rect 9413 1921 9447 1955
rect 5917 1853 5951 1887
rect 6101 1853 6135 1887
rect 6929 1853 6963 1887
rect 7113 1853 7147 1887
rect 7205 1853 7239 1887
rect 7297 1853 7331 1887
rect 8401 1853 8435 1887
rect 9505 1853 9539 1887
rect 4506 1785 4540 1819
rect 6377 1785 6411 1819
rect 6593 1785 6627 1819
rect 7665 1785 7699 1819
rect 7849 1785 7883 1819
rect 8033 1785 8067 1819
rect 9597 1785 9631 1819
rect 6745 1717 6779 1751
rect 7573 1717 7607 1751
rect 4537 1513 4571 1547
rect 4705 1513 4739 1547
rect 5825 1513 5859 1547
rect 8677 1513 8711 1547
rect 4905 1445 4939 1479
rect 6938 1445 6972 1479
rect 7205 1377 7239 1411
rect 7297 1377 7331 1411
rect 7564 1377 7598 1411
rect 4721 1173 4755 1207
<< metal1 >>
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 3694 9908 3700 9920
rect 3568 9880 3700 9908
rect 3568 9868 3574 9880
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 552 9818 10212 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 10212 9818
rect 552 9744 10212 9766
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4580 9676 6040 9704
rect 4580 9664 4586 9676
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 2682 9568 2688 9580
rect 2271 9540 2688 9568
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 2409 9503 2467 9509
rect 2409 9500 2421 9503
rect 1636 9472 2421 9500
rect 1636 9460 1642 9472
rect 2409 9469 2421 9472
rect 2455 9469 2467 9503
rect 2409 9463 2467 9469
rect 2866 9460 2872 9512
rect 2924 9500 2930 9512
rect 3237 9503 3295 9509
rect 3237 9500 3249 9503
rect 2924 9472 3249 9500
rect 2924 9460 2930 9472
rect 3237 9469 3249 9472
rect 3283 9469 3295 9503
rect 3237 9463 3295 9469
rect 3510 9460 3516 9512
rect 3568 9500 3574 9512
rect 3697 9503 3755 9509
rect 3697 9500 3709 9503
rect 3568 9472 3709 9500
rect 3568 9460 3574 9472
rect 3697 9469 3709 9472
rect 3743 9469 3755 9503
rect 5169 9503 5227 9509
rect 5169 9500 5181 9503
rect 3697 9463 3755 9469
rect 4264 9472 5181 9500
rect 4264 9444 4292 9472
rect 5169 9469 5181 9472
rect 5215 9469 5227 9503
rect 5169 9463 5227 9469
rect 5350 9460 5356 9512
rect 5408 9500 5414 9512
rect 6012 9509 6040 9676
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 8662 9704 8668 9716
rect 6604 9676 8668 9704
rect 6604 9664 6610 9676
rect 8662 9664 8668 9676
rect 8720 9664 8726 9716
rect 6178 9596 6184 9648
rect 6236 9636 6242 9648
rect 6236 9608 7328 9636
rect 6236 9596 6242 9608
rect 7006 9568 7012 9580
rect 6104 9540 7012 9568
rect 6104 9509 6132 9540
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 5629 9503 5687 9509
rect 5629 9500 5641 9503
rect 5408 9472 5641 9500
rect 5408 9460 5414 9472
rect 5629 9469 5641 9472
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 5997 9503 6055 9509
rect 5997 9469 6009 9503
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 6089 9503 6147 9509
rect 6089 9469 6101 9503
rect 6135 9469 6147 9503
rect 6089 9463 6147 9469
rect 6362 9460 6368 9512
rect 6420 9460 6426 9512
rect 7300 9509 7328 9608
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 7466 9460 7472 9512
rect 7524 9460 7530 9512
rect 8386 9460 8392 9512
rect 8444 9460 8450 9512
rect 1762 9392 1768 9444
rect 1820 9432 1826 9444
rect 1958 9435 2016 9441
rect 1958 9432 1970 9435
rect 1820 9404 1970 9432
rect 1820 9392 1826 9404
rect 1958 9401 1970 9404
rect 2004 9401 2016 9435
rect 1958 9395 2016 9401
rect 4246 9392 4252 9444
rect 4304 9392 4310 9444
rect 4924 9435 4982 9441
rect 4924 9401 4936 9435
rect 4970 9432 4982 9435
rect 7374 9432 7380 9444
rect 4970 9404 5856 9432
rect 4970 9401 4982 9404
rect 4924 9395 4982 9401
rect 845 9367 903 9373
rect 845 9364 857 9367
rect 492 9336 857 9364
rect 492 9024 520 9336
rect 845 9333 857 9336
rect 891 9333 903 9367
rect 845 9327 903 9333
rect 3050 9324 3056 9376
rect 3108 9324 3114 9376
rect 3326 9324 3332 9376
rect 3384 9364 3390 9376
rect 3421 9367 3479 9373
rect 3421 9364 3433 9367
rect 3384 9336 3433 9364
rect 3384 9324 3390 9336
rect 3421 9333 3433 9336
rect 3467 9333 3479 9367
rect 3421 9327 3479 9333
rect 3510 9324 3516 9376
rect 3568 9324 3574 9376
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3660 9336 3801 9364
rect 3660 9324 3666 9336
rect 3789 9333 3801 9336
rect 3835 9333 3847 9367
rect 3789 9327 3847 9333
rect 5442 9324 5448 9376
rect 5500 9324 5506 9376
rect 5828 9373 5856 9404
rect 6288 9404 7380 9432
rect 6288 9373 6316 9404
rect 7374 9392 7380 9404
rect 7432 9392 7438 9444
rect 7558 9392 7564 9444
rect 7616 9432 7622 9444
rect 8634 9435 8692 9441
rect 8634 9432 8646 9435
rect 7616 9404 8646 9432
rect 7616 9392 7622 9404
rect 8634 9401 8646 9404
rect 8680 9401 8692 9435
rect 8634 9395 8692 9401
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9333 5871 9367
rect 5813 9327 5871 9333
rect 6273 9367 6331 9373
rect 6273 9333 6285 9367
rect 6319 9333 6331 9367
rect 6273 9327 6331 9333
rect 7006 9324 7012 9376
rect 7064 9324 7070 9376
rect 7098 9324 7104 9376
rect 7156 9324 7162 9376
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 8113 9367 8171 9373
rect 8113 9364 8125 9367
rect 7800 9336 8125 9364
rect 7800 9324 7806 9336
rect 8113 9333 8125 9336
rect 8159 9333 8171 9367
rect 8113 9327 8171 9333
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 9769 9367 9827 9373
rect 9769 9364 9781 9367
rect 9732 9336 9781 9364
rect 9732 9324 9738 9336
rect 9769 9333 9781 9336
rect 9815 9333 9827 9367
rect 9769 9327 9827 9333
rect 552 9274 10212 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 10212 9274
rect 552 9200 10212 9222
rect 1578 9120 1584 9172
rect 1636 9120 1642 9172
rect 5629 9163 5687 9169
rect 5629 9129 5641 9163
rect 5675 9160 5687 9163
rect 6362 9160 6368 9172
rect 5675 9132 6368 9160
rect 5675 9129 5687 9132
rect 5629 9123 5687 9129
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 7193 9163 7251 9169
rect 7193 9129 7205 9163
rect 7239 9160 7251 9163
rect 7466 9160 7472 9172
rect 7239 9132 7472 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9160 9735 9163
rect 10318 9160 10324 9172
rect 9723 9132 10324 9160
rect 9723 9129 9735 9132
rect 9677 9123 9735 9129
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 2038 9052 2044 9104
rect 2096 9052 2102 9104
rect 2716 9095 2774 9101
rect 2716 9061 2728 9095
rect 2762 9092 2774 9095
rect 3510 9092 3516 9104
rect 2762 9064 3516 9092
rect 2762 9061 2774 9064
rect 2716 9055 2774 9061
rect 3510 9052 3516 9064
rect 3568 9052 3574 9104
rect 4516 9095 4574 9101
rect 4516 9061 4528 9095
rect 4562 9092 4574 9095
rect 5442 9092 5448 9104
rect 4562 9064 5448 9092
rect 4562 9061 4574 9064
rect 4516 9055 4574 9061
rect 5442 9052 5448 9064
rect 5500 9052 5506 9104
rect 6822 9092 6828 9104
rect 5828 9064 6828 9092
rect 845 9027 903 9033
rect 845 9024 857 9027
rect 492 8996 857 9024
rect 845 8993 857 8996
rect 891 8993 903 9027
rect 2056 9024 2084 9052
rect 3237 9027 3295 9033
rect 3237 9024 3249 9027
rect 2056 8996 3249 9024
rect 845 8987 903 8993
rect 3237 8993 3249 8996
rect 3283 8993 3295 9027
rect 4246 9024 4252 9036
rect 3237 8987 3295 8993
rect 3436 8996 4252 9024
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 3436 8956 3464 8996
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 5828 9033 5856 9064
rect 6822 9052 6828 9064
rect 6880 9092 6886 9104
rect 6880 9064 7328 9092
rect 6880 9052 6886 9064
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 8993 5871 9027
rect 5813 8987 5871 8993
rect 6080 9027 6138 9033
rect 6080 8993 6092 9027
rect 6126 9024 6138 9027
rect 7098 9024 7104 9036
rect 6126 8996 7104 9024
rect 6126 8993 6138 8996
rect 6080 8987 6138 8993
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 7300 9033 7328 9064
rect 7374 9052 7380 9104
rect 7432 9092 7438 9104
rect 7552 9095 7610 9101
rect 7552 9092 7564 9095
rect 7432 9064 7564 9092
rect 7432 9052 7438 9064
rect 7552 9061 7564 9064
rect 7598 9061 7610 9095
rect 7552 9055 7610 9061
rect 7285 9027 7343 9033
rect 7285 8993 7297 9027
rect 7331 8993 7343 9027
rect 7285 8987 7343 8993
rect 9122 8984 9128 9036
rect 9180 9024 9186 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 9180 8996 9505 9024
rect 9180 8984 9186 8996
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 3007 8928 3464 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3602 8916 3608 8968
rect 3660 8916 3666 8968
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 9766 8956 9772 8968
rect 9447 8928 9772 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 8757 8891 8815 8897
rect 8757 8888 8769 8891
rect 8220 8860 8769 8888
rect 1486 8780 1492 8832
rect 1544 8780 1550 8832
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 3053 8823 3111 8829
rect 3053 8820 3065 8823
rect 2832 8792 3065 8820
rect 2832 8780 2838 8792
rect 3053 8789 3065 8792
rect 3099 8789 3111 8823
rect 3053 8783 3111 8789
rect 4157 8823 4215 8829
rect 4157 8789 4169 8823
rect 4203 8820 4215 8823
rect 4890 8820 4896 8832
rect 4203 8792 4896 8820
rect 4203 8789 4215 8792
rect 4157 8783 4215 8789
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 8220 8820 8248 8860
rect 8757 8857 8769 8860
rect 8803 8857 8815 8891
rect 8757 8851 8815 8857
rect 7156 8792 8248 8820
rect 7156 8780 7162 8792
rect 8662 8780 8668 8832
rect 8720 8780 8726 8832
rect 552 8730 10212 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 10212 8730
rect 552 8656 10212 8678
rect 1489 8619 1547 8625
rect 1489 8585 1501 8619
rect 1535 8616 1547 8619
rect 1762 8616 1768 8628
rect 1535 8588 1768 8616
rect 1535 8585 1547 8588
rect 1489 8579 1547 8585
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4617 8619 4675 8625
rect 4617 8616 4629 8619
rect 4212 8588 4629 8616
rect 4212 8576 4218 8588
rect 4617 8585 4629 8588
rect 4663 8585 4675 8619
rect 4617 8579 4675 8585
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 7558 8616 7564 8628
rect 6779 8588 7564 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 9766 8576 9772 8628
rect 9824 8576 9830 8628
rect 6181 8551 6239 8557
rect 6181 8517 6193 8551
rect 6227 8548 6239 8551
rect 6270 8548 6276 8560
rect 6227 8520 6276 8548
rect 6227 8517 6239 8520
rect 6181 8511 6239 8517
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 4246 8440 4252 8492
rect 4304 8480 4310 8492
rect 4801 8483 4859 8489
rect 4801 8480 4813 8483
rect 4304 8452 4813 8480
rect 4304 8440 4310 8452
rect 4801 8449 4813 8452
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 6822 8440 6828 8492
rect 6880 8440 6886 8492
rect 382 8372 388 8424
rect 440 8412 446 8424
rect 845 8415 903 8421
rect 845 8412 857 8415
rect 440 8384 857 8412
rect 440 8372 446 8384
rect 845 8381 857 8384
rect 891 8381 903 8415
rect 845 8375 903 8381
rect 1210 8372 1216 8424
rect 1268 8412 1274 8424
rect 1305 8415 1363 8421
rect 1305 8412 1317 8415
rect 1268 8384 1317 8412
rect 1268 8372 1274 8384
rect 1305 8381 1317 8384
rect 1351 8381 1363 8415
rect 1305 8375 1363 8381
rect 1486 8372 1492 8424
rect 1544 8372 1550 8424
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8412 1639 8415
rect 2682 8412 2688 8424
rect 1627 8384 2688 8412
rect 1627 8381 1639 8384
rect 1581 8375 1639 8381
rect 2682 8372 2688 8384
rect 2740 8412 2746 8424
rect 3237 8415 3295 8421
rect 3237 8412 3249 8415
rect 2740 8384 3249 8412
rect 2740 8372 2746 8384
rect 3237 8381 3249 8384
rect 3283 8412 3295 8415
rect 4264 8412 4292 8440
rect 3283 8384 4292 8412
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 5057 8415 5115 8421
rect 5057 8412 5069 8415
rect 4948 8384 5069 8412
rect 4948 8372 4954 8384
rect 5057 8381 5069 8384
rect 5103 8381 5115 8415
rect 5057 8375 5115 8381
rect 6546 8372 6552 8424
rect 6604 8372 6610 8424
rect 6840 8412 6868 8440
rect 8386 8412 8392 8424
rect 6840 8384 8392 8412
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 1504 8344 1532 8372
rect 1826 8347 1884 8353
rect 1826 8344 1838 8347
rect 1504 8316 1838 8344
rect 1826 8313 1838 8316
rect 1872 8313 1884 8347
rect 1826 8307 1884 8313
rect 3050 8304 3056 8356
rect 3108 8344 3114 8356
rect 7098 8353 7104 8356
rect 3482 8347 3540 8353
rect 3482 8344 3494 8347
rect 3108 8316 3494 8344
rect 3108 8304 3114 8316
rect 3482 8313 3494 8316
rect 3528 8313 3540 8347
rect 7092 8344 7104 8353
rect 7059 8316 7104 8344
rect 3482 8307 3540 8313
rect 7092 8307 7104 8316
rect 7098 8304 7104 8307
rect 7156 8304 7162 8356
rect 8110 8304 8116 8356
rect 8168 8344 8174 8356
rect 8634 8347 8692 8353
rect 8634 8344 8646 8347
rect 8168 8316 8646 8344
rect 8168 8304 8174 8316
rect 8634 8313 8646 8316
rect 8680 8313 8692 8347
rect 8634 8307 8692 8313
rect 1029 8279 1087 8285
rect 1029 8245 1041 8279
rect 1075 8276 1087 8279
rect 1118 8276 1124 8288
rect 1075 8248 1124 8276
rect 1075 8245 1087 8248
rect 1029 8239 1087 8245
rect 1118 8236 1124 8248
rect 1176 8236 1182 8288
rect 2958 8236 2964 8288
rect 3016 8236 3022 8288
rect 8202 8236 8208 8288
rect 8260 8236 8266 8288
rect 552 8186 10212 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 10212 8186
rect 552 8112 10212 8134
rect 2682 8032 2688 8084
rect 2740 8032 2746 8084
rect 7006 8032 7012 8084
rect 7064 8032 7070 8084
rect 8386 8032 8392 8084
rect 8444 8072 8450 8084
rect 8665 8075 8723 8081
rect 8665 8072 8677 8075
rect 8444 8044 8677 8072
rect 8444 8032 8450 8044
rect 8665 8041 8677 8044
rect 8711 8072 8723 8075
rect 8754 8072 8760 8084
rect 8711 8044 8760 8072
rect 8711 8041 8723 8044
rect 8665 8035 8723 8041
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 3973 7939 4031 7945
rect 3973 7905 3985 7939
rect 4019 7905 4031 7939
rect 3973 7899 4031 7905
rect 6937 7939 6995 7945
rect 6937 7905 6949 7939
rect 6983 7936 6995 7939
rect 7024 7936 7052 8032
rect 6983 7908 7052 7936
rect 6983 7905 6995 7908
rect 6937 7899 6995 7905
rect 3988 7800 4016 7899
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 7156 7908 7205 7936
rect 7156 7896 7162 7908
rect 7193 7905 7205 7908
rect 7239 7905 7251 7939
rect 7193 7899 7251 7905
rect 7377 7939 7435 7945
rect 7377 7905 7389 7939
rect 7423 7905 7435 7939
rect 7377 7899 7435 7905
rect 3988 7772 6316 7800
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7732 5871 7735
rect 5994 7732 6000 7744
rect 5859 7704 6000 7732
rect 5859 7701 5871 7704
rect 5813 7695 5871 7701
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 6288 7732 6316 7772
rect 7282 7732 7288 7744
rect 6288 7704 7288 7732
rect 7282 7692 7288 7704
rect 7340 7732 7346 7744
rect 7392 7732 7420 7899
rect 8662 7896 8668 7948
rect 8720 7936 8726 7948
rect 9769 7939 9827 7945
rect 9769 7936 9781 7939
rect 8720 7908 9781 7936
rect 8720 7896 8726 7908
rect 9769 7905 9781 7908
rect 9815 7905 9827 7939
rect 9769 7899 9827 7905
rect 7340 7704 7420 7732
rect 7340 7692 7346 7704
rect 9214 7692 9220 7744
rect 9272 7692 9278 7744
rect 552 7642 10212 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 10212 7642
rect 552 7568 10212 7590
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 7156 7500 7880 7528
rect 7156 7488 7162 7500
rect 4617 7463 4675 7469
rect 4617 7429 4629 7463
rect 4663 7460 4675 7463
rect 4663 7432 5304 7460
rect 4663 7429 4675 7432
rect 4617 7423 4675 7429
rect 2682 7352 2688 7404
rect 2740 7392 2746 7404
rect 5276 7401 5304 7432
rect 7852 7401 7880 7500
rect 8110 7488 8116 7540
rect 8168 7488 8174 7540
rect 3237 7395 3295 7401
rect 3237 7392 3249 7395
rect 2740 7364 3249 7392
rect 2740 7352 2746 7364
rect 3237 7361 3249 7364
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 5261 7395 5319 7401
rect 5261 7361 5273 7395
rect 5307 7361 5319 7395
rect 5261 7355 5319 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 1118 7333 1124 7336
rect 845 7327 903 7333
rect 845 7293 857 7327
rect 891 7293 903 7327
rect 845 7287 903 7293
rect 1112 7287 1124 7333
rect 1176 7324 1182 7336
rect 1176 7296 1212 7324
rect 860 7188 888 7287
rect 1118 7284 1124 7287
rect 1176 7284 1182 7296
rect 3326 7284 3332 7336
rect 3384 7324 3390 7336
rect 3493 7327 3551 7333
rect 3493 7324 3505 7327
rect 3384 7296 3505 7324
rect 3384 7284 3390 7296
rect 3493 7293 3505 7296
rect 3539 7293 3551 7327
rect 3493 7287 3551 7293
rect 5994 7284 6000 7336
rect 6052 7284 6058 7336
rect 7581 7327 7639 7333
rect 7581 7293 7593 7327
rect 7627 7324 7639 7327
rect 7742 7324 7748 7336
rect 7627 7296 7748 7324
rect 7627 7293 7639 7296
rect 7581 7287 7639 7293
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7293 7987 7327
rect 7929 7287 7987 7293
rect 7834 7216 7840 7268
rect 7892 7256 7898 7268
rect 7944 7256 7972 7287
rect 8754 7284 8760 7336
rect 8812 7324 8818 7336
rect 9861 7327 9919 7333
rect 9861 7324 9873 7327
rect 8812 7296 9873 7324
rect 8812 7284 8818 7296
rect 9861 7293 9873 7296
rect 9907 7293 9919 7327
rect 9861 7287 9919 7293
rect 7892 7228 7972 7256
rect 7892 7216 7898 7228
rect 9490 7216 9496 7268
rect 9548 7256 9554 7268
rect 9594 7259 9652 7265
rect 9594 7256 9606 7259
rect 9548 7228 9606 7256
rect 9548 7216 9554 7228
rect 9594 7225 9606 7228
rect 9640 7225 9652 7259
rect 9594 7219 9652 7225
rect 2130 7188 2136 7200
rect 860 7160 2136 7188
rect 2130 7148 2136 7160
rect 2188 7148 2194 7200
rect 2225 7191 2283 7197
rect 2225 7157 2237 7191
rect 2271 7188 2283 7191
rect 2866 7188 2872 7200
rect 2271 7160 2872 7188
rect 2271 7157 2283 7160
rect 2225 7151 2283 7157
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 4706 7148 4712 7200
rect 4764 7148 4770 7200
rect 5994 7148 6000 7200
rect 6052 7188 6058 7200
rect 6089 7191 6147 7197
rect 6089 7188 6101 7191
rect 6052 7160 6101 7188
rect 6052 7148 6058 7160
rect 6089 7157 6101 7160
rect 6135 7157 6147 7191
rect 6089 7151 6147 7157
rect 6457 7191 6515 7197
rect 6457 7157 6469 7191
rect 6503 7188 6515 7191
rect 6546 7188 6552 7200
rect 6503 7160 6552 7188
rect 6503 7157 6515 7160
rect 6457 7151 6515 7157
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 8478 7148 8484 7200
rect 8536 7148 8542 7200
rect 552 7098 10212 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 10212 7098
rect 552 7024 10212 7046
rect 8512 6919 8570 6925
rect 8512 6885 8524 6919
rect 8558 6916 8570 6919
rect 9214 6916 9220 6928
rect 8558 6888 9220 6916
rect 8558 6885 8570 6888
rect 8512 6879 8570 6885
rect 9214 6876 9220 6888
rect 9272 6876 9278 6928
rect 1969 6851 2027 6857
rect 1969 6817 1981 6851
rect 2015 6848 2027 6851
rect 2774 6848 2780 6860
rect 2015 6820 2780 6848
rect 2015 6817 2027 6820
rect 1969 6811 2027 6817
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 2866 6808 2872 6860
rect 2924 6808 2930 6860
rect 3872 6851 3930 6857
rect 3872 6817 3884 6851
rect 3918 6848 3930 6851
rect 4706 6848 4712 6860
rect 3918 6820 4712 6848
rect 3918 6817 3930 6820
rect 3872 6811 3930 6817
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 8754 6808 8760 6860
rect 8812 6808 8818 6860
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9858 6848 9864 6860
rect 9539 6820 9864 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 2222 6740 2228 6792
rect 2280 6780 2286 6792
rect 2682 6780 2688 6792
rect 2280 6752 2688 6780
rect 2280 6740 2286 6752
rect 2682 6740 2688 6752
rect 2740 6740 2746 6792
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6749 3663 6783
rect 3605 6743 3663 6749
rect 3620 6712 3648 6743
rect 2240 6684 3648 6712
rect 845 6647 903 6653
rect 845 6644 857 6647
rect 492 6616 857 6644
rect 492 6304 520 6616
rect 845 6613 857 6616
rect 891 6613 903 6647
rect 845 6607 903 6613
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 2240 6644 2268 6684
rect 9582 6672 9588 6724
rect 9640 6712 9646 6724
rect 9677 6715 9735 6721
rect 9677 6712 9689 6715
rect 9640 6684 9689 6712
rect 9640 6672 9646 6684
rect 9677 6681 9689 6684
rect 9723 6681 9735 6715
rect 9677 6675 9735 6681
rect 1912 6616 2268 6644
rect 1912 6604 1918 6616
rect 2314 6604 2320 6656
rect 2372 6604 2378 6656
rect 4982 6604 4988 6656
rect 5040 6604 5046 6656
rect 7377 6647 7435 6653
rect 7377 6613 7389 6647
rect 7423 6644 7435 6647
rect 7742 6644 7748 6656
rect 7423 6616 7748 6644
rect 7423 6613 7435 6616
rect 7377 6607 7435 6613
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 8846 6604 8852 6656
rect 8904 6604 8910 6656
rect 552 6554 10212 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 10212 6554
rect 552 6480 10212 6502
rect 3789 6443 3847 6449
rect 3789 6409 3801 6443
rect 3835 6440 3847 6443
rect 7190 6440 7196 6452
rect 3835 6412 7196 6440
rect 3835 6409 3847 6412
rect 3789 6403 3847 6409
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 8754 6440 8760 6452
rect 7392 6412 8760 6440
rect 7392 6384 7420 6412
rect 3970 6372 3976 6384
rect 3528 6344 3976 6372
rect 3528 6313 3556 6344
rect 3970 6332 3976 6344
rect 4028 6372 4034 6384
rect 4341 6375 4399 6381
rect 4341 6372 4353 6375
rect 4028 6344 4353 6372
rect 4028 6332 4034 6344
rect 4341 6341 4353 6344
rect 4387 6341 4399 6375
rect 4341 6335 4399 6341
rect 6914 6332 6920 6384
rect 6972 6372 6978 6384
rect 7101 6375 7159 6381
rect 7101 6372 7113 6375
rect 6972 6344 7113 6372
rect 6972 6332 6978 6344
rect 7101 6341 7113 6344
rect 7147 6341 7159 6375
rect 7101 6335 7159 6341
rect 7374 6332 7380 6384
rect 7432 6332 7438 6384
rect 7745 6375 7803 6381
rect 7745 6341 7757 6375
rect 7791 6341 7803 6375
rect 7745 6335 7803 6341
rect 937 6307 995 6313
rect 937 6304 949 6307
rect 492 6276 949 6304
rect 937 6273 949 6276
rect 983 6273 995 6307
rect 937 6267 995 6273
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6304 5779 6307
rect 7392 6304 7420 6332
rect 5767 6276 7420 6304
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 2222 6236 2228 6248
rect 1719 6208 2228 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 2222 6196 2228 6208
rect 2280 6196 2286 6248
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 3016 6208 3433 6236
rect 3016 6196 3022 6208
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3421 6199 3479 6205
rect 6086 6196 6092 6248
rect 6144 6196 6150 6248
rect 6362 6196 6368 6248
rect 6420 6196 6426 6248
rect 6546 6196 6552 6248
rect 6604 6236 6610 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6604 6208 6837 6236
rect 6604 6196 6610 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 6825 6199 6883 6205
rect 6932 6208 7297 6236
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6168 1639 6171
rect 1918 6171 1976 6177
rect 1918 6168 1930 6171
rect 1627 6140 1930 6168
rect 1627 6137 1639 6140
rect 1581 6131 1639 6137
rect 1918 6137 1930 6140
rect 1964 6137 1976 6171
rect 1918 6131 1976 6137
rect 5476 6171 5534 6177
rect 5476 6137 5488 6171
rect 5522 6168 5534 6171
rect 5522 6140 5672 6168
rect 5522 6137 5534 6140
rect 5476 6131 5534 6137
rect 3053 6103 3111 6109
rect 3053 6069 3065 6103
rect 3099 6100 3111 6103
rect 3234 6100 3240 6112
rect 3099 6072 3240 6100
rect 3099 6069 3111 6072
rect 3053 6063 3111 6069
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 5644 6100 5672 6140
rect 5810 6128 5816 6180
rect 5868 6128 5874 6180
rect 6380 6168 6408 6196
rect 6641 6171 6699 6177
rect 6641 6168 6653 6171
rect 6380 6140 6653 6168
rect 6641 6137 6653 6140
rect 6687 6137 6699 6171
rect 6641 6131 6699 6137
rect 5911 6103 5969 6109
rect 5911 6100 5923 6103
rect 5644 6072 5923 6100
rect 5911 6069 5923 6072
rect 5957 6069 5969 6103
rect 5911 6063 5969 6069
rect 5997 6103 6055 6109
rect 5997 6069 6009 6103
rect 6043 6100 6055 6103
rect 6178 6100 6184 6112
rect 6043 6072 6184 6100
rect 6043 6069 6055 6072
rect 5997 6063 6055 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 6549 6103 6607 6109
rect 6549 6069 6561 6103
rect 6595 6100 6607 6103
rect 6932 6100 6960 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 7377 6239 7435 6245
rect 7377 6205 7389 6239
rect 7423 6205 7435 6239
rect 7377 6199 7435 6205
rect 7101 6171 7159 6177
rect 7101 6137 7113 6171
rect 7147 6168 7159 6171
rect 7190 6168 7196 6180
rect 7147 6140 7196 6168
rect 7147 6137 7159 6140
rect 7101 6131 7159 6137
rect 7190 6128 7196 6140
rect 7248 6128 7254 6180
rect 6595 6072 6960 6100
rect 7009 6103 7067 6109
rect 6595 6069 6607 6072
rect 6549 6063 6607 6069
rect 7009 6069 7021 6103
rect 7055 6100 7067 6103
rect 7392 6100 7420 6199
rect 7466 6196 7472 6248
rect 7524 6196 7530 6248
rect 7760 6236 7788 6335
rect 8404 6313 8432 6412
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 9858 6440 9864 6452
rect 9815 6412 9864 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 8645 6239 8703 6245
rect 8645 6236 8657 6239
rect 7760 6208 8657 6236
rect 8645 6205 8657 6208
rect 8691 6205 8703 6239
rect 8645 6199 8703 6205
rect 7650 6128 7656 6180
rect 7708 6168 7714 6180
rect 7745 6171 7803 6177
rect 7745 6168 7757 6171
rect 7708 6140 7757 6168
rect 7708 6128 7714 6140
rect 7745 6137 7757 6140
rect 7791 6137 7803 6171
rect 7745 6131 7803 6137
rect 7055 6072 7420 6100
rect 7055 6069 7067 6072
rect 7009 6063 7067 6069
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 8846 6100 8852 6112
rect 7616 6072 8852 6100
rect 7616 6060 7622 6072
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 552 6010 10212 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 10212 6010
rect 552 5936 10212 5958
rect 5537 5899 5595 5905
rect 5537 5865 5549 5899
rect 5583 5896 5595 5899
rect 5810 5896 5816 5908
rect 5583 5868 5816 5896
rect 5583 5865 5595 5868
rect 5537 5859 5595 5865
rect 5810 5856 5816 5868
rect 5868 5856 5874 5908
rect 6726 5899 6784 5905
rect 6726 5865 6738 5899
rect 6772 5896 6784 5899
rect 7650 5896 7656 5908
rect 6772 5868 7656 5896
rect 6772 5865 6784 5868
rect 6726 5859 6784 5865
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 9122 5856 9128 5908
rect 9180 5856 9186 5908
rect 9217 5899 9275 5905
rect 9217 5865 9229 5899
rect 9263 5896 9275 5899
rect 9490 5896 9496 5908
rect 9263 5868 9496 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 2124 5831 2182 5837
rect 2124 5797 2136 5831
rect 2170 5828 2182 5831
rect 2314 5828 2320 5840
rect 2170 5800 2320 5828
rect 2170 5797 2182 5800
rect 2124 5791 2182 5797
rect 2314 5788 2320 5800
rect 2372 5788 2378 5840
rect 3326 5788 3332 5840
rect 3384 5828 3390 5840
rect 3970 5828 3976 5840
rect 3384 5800 3976 5828
rect 3384 5788 3390 5800
rect 3970 5788 3976 5800
rect 4028 5828 4034 5840
rect 6457 5831 6515 5837
rect 4028 5800 4936 5828
rect 4028 5788 4034 5800
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4908 5769 4936 5800
rect 6457 5797 6469 5831
rect 6503 5828 6515 5831
rect 7285 5831 7343 5837
rect 7285 5828 7297 5831
rect 6503 5800 7297 5828
rect 6503 5797 6515 5800
rect 6457 5791 6515 5797
rect 7285 5797 7297 5800
rect 7331 5828 7343 5831
rect 7466 5828 7472 5840
rect 7331 5800 7472 5828
rect 7331 5797 7343 5800
rect 7285 5791 7343 5797
rect 7466 5788 7472 5800
rect 7524 5788 7530 5840
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4212 5732 4445 5760
rect 4212 5720 4218 5732
rect 4433 5729 4445 5732
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 4893 5763 4951 5769
rect 4893 5729 4905 5763
rect 4939 5729 4951 5763
rect 6086 5760 6092 5772
rect 4893 5723 4951 5729
rect 5644 5732 6092 5760
rect 1762 5652 1768 5704
rect 1820 5692 1826 5704
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1820 5664 1869 5692
rect 1820 5652 1826 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 4246 5652 4252 5704
rect 4304 5652 4310 5704
rect 4798 5652 4804 5704
rect 4856 5652 4862 5704
rect 5644 5636 5672 5732
rect 6086 5720 6092 5732
rect 6144 5760 6150 5772
rect 6273 5763 6331 5769
rect 6273 5760 6285 5763
rect 6144 5732 6285 5760
rect 6144 5720 6150 5732
rect 6273 5729 6285 5732
rect 6319 5760 6331 5763
rect 6549 5763 6607 5769
rect 6549 5760 6561 5763
rect 6319 5732 6561 5760
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 6549 5729 6561 5732
rect 6595 5729 6607 5763
rect 6549 5723 6607 5729
rect 6641 5763 6699 5769
rect 6641 5729 6653 5763
rect 6687 5729 6699 5763
rect 6641 5723 6699 5729
rect 6825 5763 6883 5769
rect 6825 5729 6837 5763
rect 6871 5760 6883 5763
rect 6871 5732 7144 5760
rect 6871 5729 6883 5732
rect 6825 5723 6883 5729
rect 5813 5695 5871 5701
rect 5813 5661 5825 5695
rect 5859 5661 5871 5695
rect 5813 5655 5871 5661
rect 4709 5627 4767 5633
rect 4709 5593 4721 5627
rect 4755 5624 4767 5627
rect 5626 5624 5632 5636
rect 4755 5596 5632 5624
rect 4755 5593 4767 5596
rect 4709 5587 4767 5593
rect 5626 5584 5632 5596
rect 5684 5584 5690 5636
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5556 3295 5559
rect 5828 5556 5856 5655
rect 6178 5652 6184 5704
rect 6236 5652 6242 5704
rect 6196 5624 6224 5652
rect 6656 5624 6684 5723
rect 7006 5652 7012 5704
rect 7064 5652 7070 5704
rect 7116 5692 7144 5732
rect 7190 5720 7196 5772
rect 7248 5720 7254 5772
rect 7374 5720 7380 5772
rect 7432 5760 7438 5772
rect 7745 5763 7803 5769
rect 7745 5760 7757 5763
rect 7432 5732 7757 5760
rect 7432 5720 7438 5732
rect 7745 5729 7757 5732
rect 7791 5729 7803 5763
rect 8001 5763 8059 5769
rect 8001 5760 8013 5763
rect 7745 5723 7803 5729
rect 7852 5732 8013 5760
rect 7558 5692 7564 5704
rect 7116 5664 7564 5692
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 7852 5692 7880 5732
rect 8001 5729 8013 5732
rect 8047 5729 8059 5763
rect 8001 5723 8059 5729
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 9769 5763 9827 5769
rect 9769 5760 9781 5763
rect 9732 5732 9781 5760
rect 9732 5720 9738 5732
rect 9769 5729 9781 5732
rect 9815 5729 9827 5763
rect 9769 5723 9827 5729
rect 7668 5664 7880 5692
rect 6822 5624 6828 5636
rect 6196 5596 6828 5624
rect 6822 5584 6828 5596
rect 6880 5584 6886 5636
rect 7668 5633 7696 5664
rect 7653 5627 7711 5633
rect 7653 5593 7665 5627
rect 7699 5593 7711 5627
rect 7653 5587 7711 5593
rect 3283 5528 5856 5556
rect 3283 5525 3295 5528
rect 3237 5519 3295 5525
rect 7006 5516 7012 5568
rect 7064 5556 7070 5568
rect 8386 5556 8392 5568
rect 7064 5528 8392 5556
rect 7064 5516 7070 5528
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 552 5466 10212 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 10212 5466
rect 552 5392 10212 5414
rect 8386 5312 8392 5364
rect 8444 5312 8450 5364
rect 3326 5216 3332 5228
rect 3252 5188 3332 5216
rect 3142 5108 3148 5160
rect 3200 5148 3206 5160
rect 3252 5157 3280 5188
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 5592 5188 6561 5216
rect 5592 5176 5598 5188
rect 6549 5185 6561 5188
rect 6595 5216 6607 5219
rect 7282 5216 7288 5228
rect 6595 5188 7288 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 9033 5219 9091 5225
rect 9033 5185 9045 5219
rect 9079 5216 9091 5219
rect 9122 5216 9128 5228
rect 9079 5188 9128 5216
rect 9079 5185 9091 5188
rect 9033 5179 9091 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 3237 5151 3295 5157
rect 3237 5148 3249 5151
rect 3200 5120 3249 5148
rect 3200 5108 3206 5120
rect 3237 5117 3249 5120
rect 3283 5117 3295 5151
rect 3237 5111 3295 5117
rect 3418 5108 3424 5160
rect 3476 5108 3482 5160
rect 5626 5108 5632 5160
rect 5684 5148 5690 5160
rect 6641 5151 6699 5157
rect 6641 5148 6653 5151
rect 5684 5120 6653 5148
rect 5684 5108 5690 5120
rect 6641 5117 6653 5120
rect 6687 5117 6699 5151
rect 6641 5111 6699 5117
rect 6822 5108 6828 5160
rect 6880 5108 6886 5160
rect 2682 5040 2688 5092
rect 2740 5040 2746 5092
rect 2869 5083 2927 5089
rect 2869 5049 2881 5083
rect 2915 5080 2927 5083
rect 2958 5080 2964 5092
rect 2915 5052 2964 5080
rect 2915 5049 2927 5052
rect 2869 5043 2927 5049
rect 2958 5040 2964 5052
rect 3016 5080 3022 5092
rect 3329 5083 3387 5089
rect 3329 5080 3341 5083
rect 3016 5052 3341 5080
rect 3016 5040 3022 5052
rect 3329 5049 3341 5052
rect 3375 5049 3387 5083
rect 3329 5043 3387 5049
rect 4801 5083 4859 5089
rect 4801 5049 4813 5083
rect 4847 5080 4859 5083
rect 5350 5080 5356 5092
rect 4847 5052 5356 5080
rect 4847 5049 4859 5052
rect 4801 5043 4859 5049
rect 5350 5040 5356 5052
rect 5408 5040 5414 5092
rect 7006 5040 7012 5092
rect 7064 5040 7070 5092
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2501 5015 2559 5021
rect 2501 5012 2513 5015
rect 2372 4984 2513 5012
rect 2372 4972 2378 4984
rect 2501 4981 2513 4984
rect 2547 4981 2559 5015
rect 2501 4975 2559 4981
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 6086 5012 6092 5024
rect 4764 4984 6092 5012
rect 4764 4972 4770 4984
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 552 4922 10212 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 10212 4922
rect 552 4848 10212 4870
rect 4154 4768 4160 4820
rect 4212 4768 4218 4820
rect 4706 4808 4712 4820
rect 4448 4780 4712 4808
rect 1762 4740 1768 4752
rect 952 4712 1768 4740
rect 952 4681 980 4712
rect 1762 4700 1768 4712
rect 1820 4700 1826 4752
rect 2685 4743 2743 4749
rect 2685 4709 2697 4743
rect 2731 4740 2743 4743
rect 2774 4740 2780 4752
rect 2731 4712 2780 4740
rect 2731 4709 2743 4712
rect 2685 4703 2743 4709
rect 2774 4700 2780 4712
rect 2832 4740 2838 4752
rect 3142 4740 3148 4752
rect 2832 4712 3148 4740
rect 2832 4700 2838 4712
rect 3142 4700 3148 4712
rect 3200 4700 3206 4752
rect 3326 4700 3332 4752
rect 3384 4740 3390 4752
rect 3789 4743 3847 4749
rect 3789 4740 3801 4743
rect 3384 4712 3801 4740
rect 3384 4700 3390 4712
rect 3789 4709 3801 4712
rect 3835 4709 3847 4743
rect 3789 4703 3847 4709
rect 3973 4743 4031 4749
rect 3973 4709 3985 4743
rect 4019 4740 4031 4743
rect 4062 4740 4068 4752
rect 4019 4712 4068 4740
rect 4019 4709 4031 4712
rect 3973 4703 4031 4709
rect 4062 4700 4068 4712
rect 4120 4700 4126 4752
rect 1210 4681 1216 4684
rect 937 4675 995 4681
rect 937 4641 949 4675
rect 983 4641 995 4675
rect 937 4635 995 4641
rect 1204 4635 1216 4681
rect 1210 4632 1216 4635
rect 1268 4632 1274 4684
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4641 2559 4675
rect 2501 4635 2559 4641
rect 2516 4604 2544 4635
rect 3234 4632 3240 4684
rect 3292 4632 3298 4684
rect 4448 4681 4476 4780
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 4798 4768 4804 4820
rect 4856 4808 4862 4820
rect 4893 4811 4951 4817
rect 4893 4808 4905 4811
rect 4856 4780 4905 4808
rect 4856 4768 4862 4780
rect 4893 4777 4905 4780
rect 4939 4777 4951 4811
rect 4893 4771 4951 4777
rect 5445 4811 5503 4817
rect 5445 4777 5457 4811
rect 5491 4808 5503 4811
rect 5626 4808 5632 4820
rect 5491 4780 5632 4808
rect 5491 4777 5503 4780
rect 5445 4771 5503 4777
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 6914 4768 6920 4820
rect 6972 4768 6978 4820
rect 7009 4811 7067 4817
rect 7009 4777 7021 4811
rect 7055 4808 7067 4811
rect 7377 4811 7435 4817
rect 7377 4808 7389 4811
rect 7055 4780 7389 4808
rect 7055 4777 7067 4780
rect 7009 4771 7067 4777
rect 7377 4777 7389 4780
rect 7423 4777 7435 4811
rect 7377 4771 7435 4777
rect 4522 4700 4528 4752
rect 4580 4700 4586 4752
rect 4617 4743 4675 4749
rect 4617 4709 4629 4743
rect 4663 4740 4675 4743
rect 4982 4740 4988 4752
rect 4663 4712 4988 4740
rect 4663 4709 4675 4712
rect 4617 4703 4675 4709
rect 4982 4700 4988 4712
rect 5040 4700 5046 4752
rect 5718 4700 5724 4752
rect 5776 4740 5782 4752
rect 6825 4743 6883 4749
rect 6825 4740 6837 4743
rect 5776 4712 6837 4740
rect 5776 4700 5782 4712
rect 6825 4709 6837 4712
rect 6871 4709 6883 4743
rect 6825 4703 6883 4709
rect 4798 4681 4804 4684
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4641 4307 4675
rect 4249 4635 4307 4641
rect 4397 4675 4476 4681
rect 4397 4641 4409 4675
rect 4443 4644 4476 4675
rect 4753 4675 4804 4681
rect 4753 4674 4765 4675
rect 4729 4644 4765 4674
rect 4443 4641 4455 4644
rect 4397 4635 4455 4641
rect 4753 4641 4765 4644
rect 4799 4641 4804 4675
rect 4753 4635 4804 4641
rect 3329 4607 3387 4613
rect 3329 4604 3341 4607
rect 2332 4576 3341 4604
rect 2332 4545 2360 4576
rect 3329 4573 3341 4576
rect 3375 4604 3387 4607
rect 3418 4604 3424 4616
rect 3375 4576 3424 4604
rect 3375 4573 3387 4576
rect 3329 4567 3387 4573
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 3605 4607 3663 4613
rect 3605 4573 3617 4607
rect 3651 4604 3663 4607
rect 4264 4604 4292 4635
rect 4798 4632 4804 4635
rect 4856 4632 4862 4684
rect 5504 4675 5562 4681
rect 5504 4641 5516 4675
rect 5550 4672 5562 4675
rect 5550 4641 5580 4672
rect 5504 4635 5580 4641
rect 3651 4576 4292 4604
rect 3651 4573 3663 4576
rect 3605 4567 3663 4573
rect 4890 4564 4896 4616
rect 4948 4604 4954 4616
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 4948 4576 4997 4604
rect 4948 4564 4954 4576
rect 4985 4573 4997 4576
rect 5031 4573 5043 4607
rect 4985 4567 5043 4573
rect 2317 4539 2375 4545
rect 2317 4505 2329 4539
rect 2363 4505 2375 4539
rect 2317 4499 2375 4505
rect 2866 4428 2872 4480
rect 2924 4428 2930 4480
rect 5077 4471 5135 4477
rect 5077 4437 5089 4471
rect 5123 4468 5135 4471
rect 5258 4468 5264 4480
rect 5123 4440 5264 4468
rect 5123 4437 5135 4440
rect 5077 4431 5135 4437
rect 5258 4428 5264 4440
rect 5316 4428 5322 4480
rect 5552 4468 5580 4635
rect 5810 4632 5816 4684
rect 5868 4632 5874 4684
rect 5994 4632 6000 4684
rect 6052 4632 6058 4684
rect 6086 4632 6092 4684
rect 6144 4632 6150 4684
rect 6270 4632 6276 4684
rect 6328 4672 6334 4684
rect 6365 4675 6423 4681
rect 6365 4672 6377 4675
rect 6328 4644 6377 4672
rect 6328 4632 6334 4644
rect 6365 4641 6377 4644
rect 6411 4672 6423 4675
rect 7650 4672 7656 4684
rect 6411 4644 7656 4672
rect 6411 4641 6423 4644
rect 6365 4635 6423 4641
rect 7650 4632 7656 4644
rect 7708 4632 7714 4684
rect 7742 4632 7748 4684
rect 7800 4632 7806 4684
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 9125 4675 9183 4681
rect 9125 4672 9137 4675
rect 8536 4644 9137 4672
rect 8536 4632 8542 4644
rect 9125 4641 9137 4644
rect 9171 4641 9183 4675
rect 9125 4635 9183 4641
rect 6178 4564 6184 4616
rect 6236 4564 6242 4616
rect 7466 4604 7472 4616
rect 6472 4576 7472 4604
rect 5629 4539 5687 4545
rect 5629 4505 5641 4539
rect 5675 4536 5687 4539
rect 6472 4536 6500 4576
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4604 7895 4607
rect 8202 4604 8208 4616
rect 7883 4576 8208 4604
rect 7883 4573 7895 4576
rect 7837 4567 7895 4573
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 9766 4604 9772 4616
rect 9263 4576 9772 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 5675 4508 6500 4536
rect 6549 4539 6607 4545
rect 5675 4505 5687 4508
rect 5629 4499 5687 4505
rect 6549 4505 6561 4539
rect 6595 4536 6607 4539
rect 7193 4539 7251 4545
rect 7193 4536 7205 4539
rect 6595 4508 7205 4536
rect 6595 4505 6607 4508
rect 6549 4499 6607 4505
rect 7193 4505 7205 4508
rect 7239 4505 7251 4539
rect 7193 4499 7251 4505
rect 7558 4496 7564 4548
rect 7616 4536 7622 4548
rect 8757 4539 8815 4545
rect 8757 4536 8769 4539
rect 7616 4508 8769 4536
rect 7616 4496 7622 4508
rect 8757 4505 8769 4508
rect 8803 4505 8815 4539
rect 8757 4499 8815 4505
rect 6641 4471 6699 4477
rect 6641 4468 6653 4471
rect 5552 4440 6653 4468
rect 6641 4437 6653 4440
rect 6687 4468 6699 4471
rect 6822 4468 6828 4480
rect 6687 4440 6828 4468
rect 6687 4437 6699 4440
rect 6641 4431 6699 4437
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 552 4378 10212 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 10212 4378
rect 552 4304 10212 4326
rect 2866 4224 2872 4276
rect 2924 4224 2930 4276
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 8849 4267 8907 4273
rect 8849 4264 8861 4267
rect 5868 4236 8861 4264
rect 5868 4224 5874 4236
rect 8849 4233 8861 4236
rect 8895 4233 8907 4267
rect 8849 4227 8907 4233
rect 5626 4156 5632 4208
rect 5684 4196 5690 4208
rect 7653 4199 7711 4205
rect 7653 4196 7665 4199
rect 5684 4168 7665 4196
rect 5684 4156 5690 4168
rect 7653 4165 7665 4168
rect 7699 4165 7711 4199
rect 7653 4159 7711 4165
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4128 3387 4131
rect 4246 4128 4252 4140
rect 3375 4100 4252 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 7837 4131 7895 4137
rect 7837 4128 7849 4131
rect 5040 4100 5856 4128
rect 5040 4088 5046 4100
rect 1213 4063 1271 4069
rect 1213 4029 1225 4063
rect 1259 4060 1271 4063
rect 1762 4060 1768 4072
rect 1259 4032 1768 4060
rect 1259 4029 1271 4032
rect 1213 4023 1271 4029
rect 1762 4020 1768 4032
rect 1820 4060 1826 4072
rect 1820 4032 3188 4060
rect 1820 4020 1826 4032
rect 1480 3995 1538 4001
rect 1480 3961 1492 3995
rect 1526 3992 1538 3995
rect 2130 3992 2136 4004
rect 1526 3964 2136 3992
rect 1526 3961 1538 3964
rect 1480 3955 1538 3961
rect 2130 3952 2136 3964
rect 2188 3952 2194 4004
rect 2853 3995 2911 4001
rect 2240 3964 2728 3992
rect 1210 3884 1216 3936
rect 1268 3924 1274 3936
rect 2240 3924 2268 3964
rect 1268 3896 2268 3924
rect 1268 3884 1274 3896
rect 2590 3884 2596 3936
rect 2648 3884 2654 3936
rect 2700 3933 2728 3964
rect 2853 3961 2865 3995
rect 2899 3992 2911 3995
rect 2958 3992 2964 4004
rect 2899 3964 2964 3992
rect 2899 3961 2911 3964
rect 2853 3955 2911 3961
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 3053 3995 3111 4001
rect 3053 3961 3065 3995
rect 3099 3961 3111 3995
rect 3160 3992 3188 4032
rect 3234 4020 3240 4072
rect 3292 4020 3298 4072
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4060 3479 4063
rect 4062 4060 4068 4072
rect 3467 4032 4068 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 5261 4063 5319 4069
rect 5261 4029 5273 4063
rect 5307 4060 5319 4063
rect 5534 4060 5540 4072
rect 5307 4032 5540 4060
rect 5307 4029 5319 4032
rect 5261 4023 5319 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 5718 4060 5724 4072
rect 5675 4032 5724 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 5828 4069 5856 4100
rect 6196 4100 7849 4128
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4029 5871 4063
rect 5813 4023 5871 4029
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4029 6055 4063
rect 5997 4023 6055 4029
rect 3160 3964 4016 3992
rect 3053 3955 3111 3961
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3893 2743 3927
rect 3068 3924 3096 3955
rect 3878 3924 3884 3936
rect 3068 3896 3884 3924
rect 2685 3887 2743 3893
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 3988 3933 4016 3964
rect 4154 3952 4160 4004
rect 4212 3992 4218 4004
rect 4798 3992 4804 4004
rect 4212 3964 4804 3992
rect 4212 3952 4218 3964
rect 4798 3952 4804 3964
rect 4856 3992 4862 4004
rect 6012 3992 6040 4023
rect 6086 4020 6092 4072
rect 6144 4020 6150 4072
rect 6196 4069 6224 4100
rect 7837 4097 7849 4100
rect 7883 4097 7895 4131
rect 7837 4091 7895 4097
rect 8018 4088 8024 4140
rect 8076 4128 8082 4140
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8076 4100 9045 4128
rect 8076 4088 8082 4100
rect 9033 4097 9045 4100
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 6181 4063 6239 4069
rect 6181 4029 6193 4063
rect 6227 4029 6239 4063
rect 6181 4023 6239 4029
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 6365 4063 6423 4069
rect 6365 4060 6377 4063
rect 6328 4032 6377 4060
rect 6328 4020 6334 4032
rect 6365 4029 6377 4032
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 6454 4020 6460 4072
rect 6512 4020 6518 4072
rect 6546 4020 6552 4072
rect 6604 4060 6610 4072
rect 7009 4063 7067 4069
rect 7009 4060 7021 4063
rect 6604 4032 7021 4060
rect 6604 4020 6610 4032
rect 7009 4029 7021 4032
rect 7055 4029 7067 4063
rect 7009 4023 7067 4029
rect 7190 4020 7196 4072
rect 7248 4020 7254 4072
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4060 7343 4063
rect 7374 4060 7380 4072
rect 7331 4032 7380 4060
rect 7331 4029 7343 4032
rect 7285 4023 7343 4029
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 7466 4020 7472 4072
rect 7524 4020 7530 4072
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 7745 4063 7803 4069
rect 7745 4060 7757 4063
rect 7708 4032 7757 4060
rect 7708 4020 7714 4032
rect 7745 4029 7757 4032
rect 7791 4029 7803 4063
rect 7745 4023 7803 4029
rect 8110 4020 8116 4072
rect 8168 4060 8174 4072
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8168 4032 9137 4060
rect 8168 4020 8174 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 4856 3964 6040 3992
rect 4856 3952 4862 3964
rect 3973 3927 4031 3933
rect 3973 3893 3985 3927
rect 4019 3924 4031 3927
rect 4246 3924 4252 3936
rect 4019 3896 4252 3924
rect 4019 3893 4031 3896
rect 3973 3887 4031 3893
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 7558 3924 7564 3936
rect 6328 3896 7564 3924
rect 6328 3884 6334 3896
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 552 3834 10212 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 10212 3834
rect 552 3760 10212 3782
rect 2041 3723 2099 3729
rect 2041 3689 2053 3723
rect 2087 3720 2099 3723
rect 2291 3723 2349 3729
rect 2291 3720 2303 3723
rect 2087 3692 2303 3720
rect 2087 3689 2099 3692
rect 2041 3683 2099 3689
rect 2291 3689 2303 3692
rect 2337 3689 2349 3723
rect 2958 3720 2964 3732
rect 2291 3683 2349 3689
rect 2424 3692 2964 3720
rect 2424 3652 2452 3692
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3145 3723 3203 3729
rect 3145 3689 3157 3723
rect 3191 3720 3203 3723
rect 3326 3720 3332 3732
rect 3191 3692 3332 3720
rect 3191 3689 3203 3692
rect 3145 3683 3203 3689
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 3418 3680 3424 3732
rect 3476 3680 3482 3732
rect 3789 3723 3847 3729
rect 3789 3689 3801 3723
rect 3835 3720 3847 3723
rect 4890 3720 4896 3732
rect 3835 3692 4896 3720
rect 3835 3689 3847 3692
rect 3789 3683 3847 3689
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 5905 3723 5963 3729
rect 5905 3689 5917 3723
rect 5951 3720 5963 3723
rect 6178 3720 6184 3732
rect 5951 3692 6184 3720
rect 5951 3689 5963 3692
rect 5905 3683 5963 3689
rect 6178 3680 6184 3692
rect 6236 3720 6242 3732
rect 7190 3720 7196 3732
rect 6236 3692 7196 3720
rect 6236 3680 6242 3692
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 7282 3680 7288 3732
rect 7340 3680 7346 3732
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 8754 3720 8760 3732
rect 8352 3692 8760 3720
rect 8352 3680 8358 3692
rect 8754 3680 8760 3692
rect 8812 3720 8818 3732
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 8812 3692 8953 3720
rect 8812 3680 8818 3692
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 8941 3683 8999 3689
rect 1872 3624 2452 3652
rect 2501 3655 2559 3661
rect 1872 3593 1900 3624
rect 2501 3621 2513 3655
rect 2547 3621 2559 3655
rect 3513 3655 3571 3661
rect 3513 3652 3525 3655
rect 2501 3615 2559 3621
rect 2976 3624 3525 3652
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 2038 3544 2044 3596
rect 2096 3544 2102 3596
rect 2516 3516 2544 3615
rect 2590 3544 2596 3596
rect 2648 3584 2654 3596
rect 2976 3593 3004 3624
rect 3513 3621 3525 3624
rect 3559 3652 3571 3655
rect 3559 3624 3924 3652
rect 3559 3621 3571 3624
rect 3513 3615 3571 3621
rect 2961 3587 3019 3593
rect 2961 3584 2973 3587
rect 2648 3556 2973 3584
rect 2648 3544 2654 3556
rect 2961 3553 2973 3556
rect 3007 3553 3019 3587
rect 2961 3547 3019 3553
rect 3050 3544 3056 3596
rect 3108 3584 3114 3596
rect 3234 3584 3240 3596
rect 3108 3556 3240 3584
rect 3108 3544 3114 3556
rect 3234 3544 3240 3556
rect 3292 3584 3298 3596
rect 3896 3593 3924 3624
rect 3970 3612 3976 3664
rect 4028 3652 4034 3664
rect 4154 3652 4160 3664
rect 4028 3624 4160 3652
rect 4028 3612 4034 3624
rect 4154 3612 4160 3624
rect 4212 3612 4218 3664
rect 4516 3655 4574 3661
rect 4516 3621 4528 3655
rect 4562 3652 4574 3655
rect 5626 3652 5632 3664
rect 4562 3624 5632 3652
rect 4562 3621 4574 3624
rect 4516 3615 4574 3621
rect 5626 3612 5632 3624
rect 5684 3612 5690 3664
rect 7300 3652 7328 3680
rect 7653 3655 7711 3661
rect 7653 3652 7665 3655
rect 7300 3624 7665 3652
rect 7653 3621 7665 3624
rect 7699 3621 7711 3655
rect 7653 3615 7711 3621
rect 3605 3587 3663 3593
rect 3605 3584 3617 3587
rect 3292 3556 3617 3584
rect 3292 3544 3298 3556
rect 3605 3553 3617 3556
rect 3651 3553 3663 3587
rect 3605 3547 3663 3553
rect 3881 3587 3939 3593
rect 3881 3553 3893 3587
rect 3927 3553 3939 3587
rect 3881 3547 3939 3553
rect 5997 3587 6055 3593
rect 5997 3553 6009 3587
rect 6043 3584 6055 3587
rect 6454 3584 6460 3596
rect 6043 3556 6460 3584
rect 6043 3553 6055 3556
rect 5997 3547 6055 3553
rect 2685 3519 2743 3525
rect 2516 3488 2636 3516
rect 2130 3408 2136 3460
rect 2188 3408 2194 3460
rect 2314 3340 2320 3392
rect 2372 3340 2378 3392
rect 2608 3380 2636 3488
rect 2685 3485 2697 3519
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 2700 3448 2728 3479
rect 2774 3476 2780 3528
rect 2832 3476 2838 3528
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3516 2927 3519
rect 3418 3516 3424 3528
rect 2915 3488 3424 3516
rect 2915 3485 2927 3488
rect 2869 3479 2927 3485
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 3510 3476 3516 3528
rect 3568 3516 3574 3528
rect 3620 3516 3648 3547
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 7006 3584 7012 3596
rect 6963 3556 7012 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 7098 3544 7104 3596
rect 7156 3544 7162 3596
rect 7193 3587 7251 3593
rect 7193 3553 7205 3587
rect 7239 3553 7251 3587
rect 7193 3547 7251 3553
rect 3568 3488 3648 3516
rect 3568 3476 3574 3488
rect 4246 3476 4252 3528
rect 4304 3476 4310 3528
rect 7208 3516 7236 3547
rect 7282 3544 7288 3596
rect 7340 3544 7346 3596
rect 8386 3516 8392 3528
rect 7208 3488 8392 3516
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 3050 3448 3056 3460
rect 2700 3420 3056 3448
rect 3050 3408 3056 3420
rect 3108 3408 3114 3460
rect 3234 3408 3240 3460
rect 3292 3408 3298 3460
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 5629 3451 5687 3457
rect 5629 3448 5641 3451
rect 5316 3420 5641 3448
rect 5316 3408 5322 3420
rect 5629 3417 5641 3420
rect 5675 3448 5687 3451
rect 6086 3448 6092 3460
rect 5675 3420 6092 3448
rect 5675 3417 5687 3420
rect 5629 3411 5687 3417
rect 6086 3408 6092 3420
rect 6144 3408 6150 3460
rect 2774 3380 2780 3392
rect 2608 3352 2780 3380
rect 2774 3340 2780 3352
rect 2832 3340 2838 3392
rect 7561 3383 7619 3389
rect 7561 3349 7573 3383
rect 7607 3380 7619 3383
rect 8478 3380 8484 3392
rect 7607 3352 8484 3380
rect 7607 3349 7619 3352
rect 7561 3343 7619 3349
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 552 3290 10212 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 10212 3290
rect 552 3216 10212 3238
rect 3510 3136 3516 3188
rect 3568 3176 3574 3188
rect 4617 3179 4675 3185
rect 4617 3176 4629 3179
rect 3568 3148 4629 3176
rect 3568 3136 3574 3148
rect 4617 3145 4629 3148
rect 4663 3145 4675 3179
rect 4617 3139 4675 3145
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 5074 3176 5080 3188
rect 4764 3148 5080 3176
rect 4764 3136 4770 3148
rect 5074 3136 5080 3148
rect 5132 3176 5138 3188
rect 5445 3179 5503 3185
rect 5445 3176 5457 3179
rect 5132 3148 5457 3176
rect 5132 3136 5138 3148
rect 5445 3145 5457 3148
rect 5491 3145 5503 3179
rect 5445 3139 5503 3145
rect 7098 3136 7104 3188
rect 7156 3176 7162 3188
rect 7653 3179 7711 3185
rect 7653 3176 7665 3179
rect 7156 3148 7665 3176
rect 7156 3136 7162 3148
rect 7653 3145 7665 3148
rect 7699 3145 7711 3179
rect 7653 3139 7711 3145
rect 7742 3136 7748 3188
rect 7800 3176 7806 3188
rect 8018 3176 8024 3188
rect 7800 3148 8024 3176
rect 7800 3136 7806 3148
rect 8018 3136 8024 3148
rect 8076 3176 8082 3188
rect 9490 3176 9496 3188
rect 8076 3148 9496 3176
rect 8076 3136 8082 3148
rect 9490 3136 9496 3148
rect 9548 3136 9554 3188
rect 9766 3136 9772 3188
rect 9824 3136 9830 3188
rect 4798 3068 4804 3120
rect 4856 3108 4862 3120
rect 7374 3108 7380 3120
rect 4856 3080 7380 3108
rect 4856 3068 4862 3080
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 7282 3000 7288 3052
rect 7340 3040 7346 3052
rect 7340 3012 7880 3040
rect 7340 3000 7346 3012
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2972 3295 2975
rect 4246 2972 4252 2984
rect 3283 2944 4252 2972
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 4246 2932 4252 2944
rect 4304 2932 4310 2984
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2972 4767 2975
rect 4890 2972 4896 2984
rect 4755 2944 4896 2972
rect 4755 2941 4767 2944
rect 4709 2935 4767 2941
rect 4890 2932 4896 2944
rect 4948 2972 4954 2984
rect 5166 2972 5172 2984
rect 4948 2944 5172 2972
rect 4948 2932 4954 2944
rect 5166 2932 5172 2944
rect 5224 2972 5230 2984
rect 7576 2981 7604 3012
rect 7561 2975 7619 2981
rect 5224 2944 5488 2972
rect 5224 2932 5230 2944
rect 3510 2913 3516 2916
rect 3504 2867 3516 2913
rect 3510 2864 3516 2867
rect 3568 2864 3574 2916
rect 4982 2864 4988 2916
rect 5040 2904 5046 2916
rect 5258 2904 5264 2916
rect 5040 2876 5264 2904
rect 5040 2864 5046 2876
rect 5258 2864 5264 2876
rect 5316 2864 5322 2916
rect 5460 2913 5488 2944
rect 7561 2941 7573 2975
rect 7607 2941 7619 2975
rect 7561 2935 7619 2941
rect 7745 2975 7803 2981
rect 7745 2941 7757 2975
rect 7791 2941 7803 2975
rect 7852 2972 7880 3012
rect 8294 3000 8300 3052
rect 8352 3040 8358 3052
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 8352 3012 8401 3040
rect 8352 3000 8358 3012
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 7852 2944 8340 2972
rect 7745 2935 7803 2941
rect 5460 2907 5519 2913
rect 5460 2876 5473 2907
rect 5461 2873 5473 2876
rect 5507 2873 5519 2907
rect 7760 2904 7788 2935
rect 7760 2876 8156 2904
rect 5461 2867 5519 2873
rect 5626 2796 5632 2848
rect 5684 2796 5690 2848
rect 7852 2845 7880 2876
rect 8018 2845 8024 2848
rect 7837 2839 7895 2845
rect 7837 2805 7849 2839
rect 7883 2805 7895 2839
rect 7837 2799 7895 2805
rect 8005 2839 8024 2845
rect 8005 2805 8017 2839
rect 8005 2799 8024 2805
rect 8018 2796 8024 2799
rect 8076 2796 8082 2848
rect 8128 2836 8156 2876
rect 8202 2864 8208 2916
rect 8260 2864 8266 2916
rect 8312 2904 8340 2944
rect 8478 2932 8484 2984
rect 8536 2972 8542 2984
rect 8645 2975 8703 2981
rect 8645 2972 8657 2975
rect 8536 2944 8657 2972
rect 8536 2932 8542 2944
rect 8645 2941 8657 2944
rect 8691 2941 8703 2975
rect 8645 2935 8703 2941
rect 8754 2904 8760 2916
rect 8312 2876 8760 2904
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 8386 2836 8392 2848
rect 8128 2808 8392 2836
rect 8386 2796 8392 2808
rect 8444 2796 8450 2848
rect 552 2746 10212 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 10212 2746
rect 552 2672 10212 2694
rect 3510 2592 3516 2644
rect 3568 2592 3574 2644
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 5261 2635 5319 2641
rect 5261 2632 5273 2635
rect 5040 2604 5273 2632
rect 5040 2592 5046 2604
rect 5261 2601 5273 2604
rect 5307 2632 5319 2635
rect 5307 2604 5948 2632
rect 5307 2601 5319 2604
rect 5261 2595 5319 2601
rect 3142 2524 3148 2576
rect 3200 2564 3206 2576
rect 3665 2567 3723 2573
rect 3665 2564 3677 2567
rect 3200 2536 3677 2564
rect 3200 2524 3206 2536
rect 3665 2533 3677 2536
rect 3711 2533 3723 2567
rect 3665 2527 3723 2533
rect 3881 2567 3939 2573
rect 3881 2533 3893 2567
rect 3927 2564 3939 2567
rect 4062 2564 4068 2576
rect 3927 2536 4068 2564
rect 3927 2533 3939 2536
rect 3881 2527 3939 2533
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 3896 2496 3924 2527
rect 4062 2524 4068 2536
rect 4120 2524 4126 2576
rect 5920 2573 5948 2604
rect 6086 2592 6092 2644
rect 6144 2632 6150 2644
rect 6181 2635 6239 2641
rect 6181 2632 6193 2635
rect 6144 2604 6193 2632
rect 6144 2592 6150 2604
rect 6181 2601 6193 2604
rect 6227 2632 6239 2635
rect 6362 2632 6368 2644
rect 6227 2604 6368 2632
rect 6227 2601 6239 2604
rect 6181 2595 6239 2601
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 7469 2635 7527 2641
rect 7064 2604 7144 2632
rect 7064 2592 7070 2604
rect 7116 2573 7144 2604
rect 7469 2601 7481 2635
rect 7515 2632 7527 2635
rect 7515 2604 8248 2632
rect 7515 2601 7527 2604
rect 7469 2595 7527 2601
rect 5905 2567 5963 2573
rect 5092 2536 5764 2564
rect 5092 2505 5120 2536
rect 2832 2468 3924 2496
rect 5077 2499 5135 2505
rect 2832 2456 2838 2468
rect 5077 2465 5089 2499
rect 5123 2465 5135 2499
rect 5077 2459 5135 2465
rect 5092 2428 5120 2459
rect 5166 2456 5172 2508
rect 5224 2496 5230 2508
rect 5353 2499 5411 2505
rect 5353 2496 5365 2499
rect 5224 2468 5365 2496
rect 5224 2456 5230 2468
rect 5353 2465 5365 2468
rect 5399 2465 5411 2499
rect 5353 2459 5411 2465
rect 5258 2428 5264 2440
rect 5092 2400 5264 2428
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5368 2428 5396 2459
rect 5626 2456 5632 2508
rect 5684 2456 5690 2508
rect 5736 2496 5764 2536
rect 5905 2533 5917 2567
rect 5951 2533 5963 2567
rect 5905 2527 5963 2533
rect 7101 2567 7159 2573
rect 7101 2533 7113 2567
rect 7147 2533 7159 2567
rect 7101 2527 7159 2533
rect 7317 2567 7375 2573
rect 7317 2533 7329 2567
rect 7363 2564 7375 2567
rect 7834 2564 7840 2576
rect 7363 2536 7840 2564
rect 7363 2533 7375 2536
rect 7317 2527 7375 2533
rect 7834 2524 7840 2536
rect 7892 2524 7898 2576
rect 7926 2524 7932 2576
rect 7984 2524 7990 2576
rect 8220 2564 8248 2604
rect 9490 2592 9496 2644
rect 9548 2592 9554 2644
rect 8380 2567 8438 2573
rect 8380 2564 8392 2567
rect 8220 2536 8392 2564
rect 8380 2533 8392 2536
rect 8426 2533 8438 2567
rect 8380 2527 8438 2533
rect 6089 2499 6147 2505
rect 6089 2496 6101 2499
rect 5736 2468 6101 2496
rect 6089 2465 6101 2468
rect 6135 2465 6147 2499
rect 6089 2459 6147 2465
rect 6273 2499 6331 2505
rect 6273 2465 6285 2499
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 6457 2499 6515 2505
rect 6457 2465 6469 2499
rect 6503 2496 6515 2499
rect 7009 2499 7067 2505
rect 7009 2496 7021 2499
rect 6503 2468 7021 2496
rect 6503 2465 6515 2468
rect 6457 2459 6515 2465
rect 7009 2465 7021 2468
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 6288 2428 6316 2459
rect 5368 2400 6316 2428
rect 7024 2428 7052 2459
rect 7742 2456 7748 2508
rect 7800 2456 7806 2508
rect 8018 2456 8024 2508
rect 8076 2456 8082 2508
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8202 2496 8208 2508
rect 8159 2468 8208 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 8036 2428 8064 2456
rect 7024 2400 8064 2428
rect 4798 2360 4804 2372
rect 3712 2332 4804 2360
rect 3712 2301 3740 2332
rect 4798 2320 4804 2332
rect 4856 2320 4862 2372
rect 7561 2363 7619 2369
rect 7561 2360 7573 2363
rect 7300 2332 7573 2360
rect 3697 2295 3755 2301
rect 3697 2261 3709 2295
rect 3743 2261 3755 2295
rect 3697 2255 3755 2261
rect 4706 2252 4712 2304
rect 4764 2292 4770 2304
rect 4893 2295 4951 2301
rect 4893 2292 4905 2295
rect 4764 2264 4905 2292
rect 4764 2252 4770 2264
rect 4893 2261 4905 2264
rect 4939 2261 4951 2295
rect 4893 2255 4951 2261
rect 5534 2252 5540 2304
rect 5592 2252 5598 2304
rect 6917 2295 6975 2301
rect 6917 2261 6929 2295
rect 6963 2292 6975 2295
rect 7006 2292 7012 2304
rect 6963 2264 7012 2292
rect 6963 2261 6975 2264
rect 6917 2255 6975 2261
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 7300 2301 7328 2332
rect 7561 2329 7573 2332
rect 7607 2329 7619 2363
rect 7561 2323 7619 2329
rect 7285 2295 7343 2301
rect 7285 2261 7297 2295
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 552 2202 10212 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 10212 2202
rect 552 2128 10212 2150
rect 5258 2048 5264 2100
rect 5316 2088 5322 2100
rect 5629 2091 5687 2097
rect 5629 2088 5641 2091
rect 5316 2060 5641 2088
rect 5316 2048 5322 2060
rect 5629 2057 5641 2060
rect 5675 2057 5687 2091
rect 5629 2051 5687 2057
rect 6273 2091 6331 2097
rect 6273 2057 6285 2091
rect 6319 2088 6331 2091
rect 6549 2091 6607 2097
rect 6549 2088 6561 2091
rect 6319 2060 6561 2088
rect 6319 2057 6331 2060
rect 6273 2051 6331 2057
rect 6549 2057 6561 2060
rect 6595 2057 6607 2091
rect 6549 2051 6607 2057
rect 7834 2048 7840 2100
rect 7892 2088 7898 2100
rect 8481 2091 8539 2097
rect 8481 2088 8493 2091
rect 7892 2060 8493 2088
rect 7892 2048 7898 2060
rect 8481 2057 8493 2060
rect 8527 2057 8539 2091
rect 8481 2051 8539 2057
rect 8754 2048 8760 2100
rect 8812 2048 8818 2100
rect 6914 2020 6920 2032
rect 6380 1992 6920 2020
rect 4246 1912 4252 1964
rect 4304 1912 4310 1964
rect 5626 1844 5632 1896
rect 5684 1884 5690 1896
rect 5905 1887 5963 1893
rect 5905 1884 5917 1887
rect 5684 1856 5917 1884
rect 5684 1844 5690 1856
rect 5905 1853 5917 1856
rect 5951 1853 5963 1887
rect 5905 1847 5963 1853
rect 6086 1844 6092 1896
rect 6144 1844 6150 1896
rect 4246 1776 4252 1828
rect 4304 1816 4310 1828
rect 6380 1825 6408 1992
rect 6914 1980 6920 1992
rect 6972 1980 6978 2032
rect 7006 1952 7012 1964
rect 6748 1924 7012 1952
rect 4494 1819 4552 1825
rect 4494 1816 4506 1819
rect 4304 1788 4506 1816
rect 4304 1776 4310 1788
rect 4494 1785 4506 1788
rect 4540 1785 4552 1819
rect 4494 1779 4552 1785
rect 6365 1819 6423 1825
rect 6365 1785 6377 1819
rect 6411 1785 6423 1819
rect 6365 1779 6423 1785
rect 6581 1819 6639 1825
rect 6581 1785 6593 1819
rect 6627 1816 6639 1819
rect 6748 1816 6776 1924
rect 7006 1912 7012 1924
rect 7064 1952 7070 1964
rect 7064 1924 7236 1952
rect 7064 1912 7070 1924
rect 6914 1844 6920 1896
rect 6972 1844 6978 1896
rect 7208 1893 7236 1924
rect 7926 1912 7932 1964
rect 7984 1952 7990 1964
rect 9401 1955 9459 1961
rect 7984 1924 8524 1952
rect 7984 1912 7990 1924
rect 7101 1887 7159 1893
rect 7101 1853 7113 1887
rect 7147 1853 7159 1887
rect 7101 1847 7159 1853
rect 7193 1887 7251 1893
rect 7193 1853 7205 1887
rect 7239 1853 7251 1887
rect 7193 1847 7251 1853
rect 7285 1887 7343 1893
rect 7285 1853 7297 1887
rect 7331 1884 7343 1887
rect 7331 1856 8340 1884
rect 7331 1853 7343 1856
rect 7285 1847 7343 1853
rect 6627 1788 6776 1816
rect 7116 1816 7144 1847
rect 7653 1819 7711 1825
rect 7653 1816 7665 1819
rect 7116 1788 7665 1816
rect 6627 1785 6639 1788
rect 6581 1779 6639 1785
rect 7653 1785 7665 1788
rect 7699 1785 7711 1819
rect 7653 1779 7711 1785
rect 7837 1819 7895 1825
rect 7837 1785 7849 1819
rect 7883 1816 7895 1819
rect 7926 1816 7932 1828
rect 7883 1788 7932 1816
rect 7883 1785 7895 1788
rect 7837 1779 7895 1785
rect 7926 1776 7932 1788
rect 7984 1776 7990 1828
rect 8018 1776 8024 1828
rect 8076 1776 8082 1828
rect 8312 1816 8340 1856
rect 8386 1844 8392 1896
rect 8444 1844 8450 1896
rect 8496 1884 8524 1924
rect 9401 1921 9413 1955
rect 9447 1952 9459 1955
rect 9766 1952 9772 1964
rect 9447 1924 9772 1952
rect 9447 1921 9459 1924
rect 9401 1915 9459 1921
rect 9766 1912 9772 1924
rect 9824 1912 9830 1964
rect 9493 1887 9551 1893
rect 9493 1884 9505 1887
rect 8496 1856 9505 1884
rect 9493 1853 9505 1856
rect 9539 1853 9551 1887
rect 9493 1847 9551 1853
rect 9585 1819 9643 1825
rect 9585 1816 9597 1819
rect 8312 1788 9597 1816
rect 9585 1785 9597 1788
rect 9631 1785 9643 1819
rect 9585 1779 9643 1785
rect 6730 1708 6736 1760
rect 6788 1708 6794 1760
rect 7558 1708 7564 1760
rect 7616 1708 7622 1760
rect 552 1658 10212 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 10212 1658
rect 552 1584 10212 1606
rect 4246 1504 4252 1556
rect 4304 1544 4310 1556
rect 4706 1553 4712 1556
rect 4525 1547 4583 1553
rect 4525 1544 4537 1547
rect 4304 1516 4537 1544
rect 4304 1504 4310 1516
rect 4525 1513 4537 1516
rect 4571 1513 4583 1547
rect 4525 1507 4583 1513
rect 4693 1547 4712 1553
rect 4693 1513 4705 1547
rect 4693 1507 4712 1513
rect 4706 1504 4712 1507
rect 4764 1504 4770 1556
rect 5813 1547 5871 1553
rect 5813 1513 5825 1547
rect 5859 1544 5871 1547
rect 6086 1544 6092 1556
rect 5859 1516 6092 1544
rect 5859 1513 5871 1516
rect 5813 1507 5871 1513
rect 6086 1504 6092 1516
rect 6144 1504 6150 1556
rect 6822 1544 6828 1556
rect 6196 1516 6828 1544
rect 4062 1436 4068 1488
rect 4120 1476 4126 1488
rect 4893 1479 4951 1485
rect 4893 1476 4905 1479
rect 4120 1448 4905 1476
rect 4120 1436 4126 1448
rect 4893 1445 4905 1448
rect 4939 1476 4951 1479
rect 6196 1476 6224 1516
rect 6822 1504 6828 1516
rect 6880 1504 6886 1556
rect 7926 1504 7932 1556
rect 7984 1544 7990 1556
rect 8665 1547 8723 1553
rect 8665 1544 8677 1547
rect 7984 1516 8677 1544
rect 7984 1504 7990 1516
rect 8665 1513 8677 1516
rect 8711 1513 8723 1547
rect 8665 1507 8723 1513
rect 4939 1448 6224 1476
rect 4939 1445 4951 1448
rect 4893 1439 4951 1445
rect 6730 1436 6736 1488
rect 6788 1476 6794 1488
rect 6926 1479 6984 1485
rect 6926 1476 6938 1479
rect 6788 1448 6938 1476
rect 6788 1436 6794 1448
rect 6926 1445 6938 1448
rect 6972 1445 6984 1479
rect 8294 1476 8300 1488
rect 6926 1439 6984 1445
rect 7300 1448 8300 1476
rect 7300 1417 7328 1448
rect 8294 1436 8300 1448
rect 8352 1436 8358 1488
rect 7558 1417 7564 1420
rect 7193 1411 7251 1417
rect 7193 1377 7205 1411
rect 7239 1408 7251 1411
rect 7285 1411 7343 1417
rect 7285 1408 7297 1411
rect 7239 1380 7297 1408
rect 7239 1377 7251 1380
rect 7193 1371 7251 1377
rect 7285 1377 7297 1380
rect 7331 1377 7343 1411
rect 7552 1408 7564 1417
rect 7519 1380 7564 1408
rect 7285 1371 7343 1377
rect 7552 1371 7564 1380
rect 7558 1368 7564 1371
rect 7616 1368 7622 1420
rect 4709 1207 4767 1213
rect 4709 1173 4721 1207
rect 4755 1204 4767 1207
rect 5534 1204 5540 1216
rect 4755 1176 5540 1204
rect 4755 1173 4767 1176
rect 4709 1167 4767 1173
rect 5534 1164 5540 1176
rect 5592 1164 5598 1216
rect 552 1114 10212 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 10212 1114
rect 552 1040 10212 1062
rect 552 570 10212 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 10212 570
rect 552 496 10212 518
<< via1 >>
rect 3516 9868 3568 9920
rect 3700 9868 3752 9920
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 4528 9664 4580 9716
rect 2688 9528 2740 9580
rect 1584 9460 1636 9512
rect 2872 9460 2924 9512
rect 3516 9460 3568 9512
rect 5356 9460 5408 9512
rect 6552 9664 6604 9716
rect 8668 9664 8720 9716
rect 6184 9596 6236 9648
rect 7012 9528 7064 9580
rect 6368 9503 6420 9512
rect 6368 9469 6377 9503
rect 6377 9469 6411 9503
rect 6411 9469 6420 9503
rect 6368 9460 6420 9469
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 1768 9392 1820 9444
rect 4252 9392 4304 9444
rect 3056 9367 3108 9376
rect 3056 9333 3065 9367
rect 3065 9333 3099 9367
rect 3099 9333 3108 9367
rect 3056 9324 3108 9333
rect 3332 9324 3384 9376
rect 3516 9367 3568 9376
rect 3516 9333 3525 9367
rect 3525 9333 3559 9367
rect 3559 9333 3568 9367
rect 3516 9324 3568 9333
rect 3608 9324 3660 9376
rect 5448 9367 5500 9376
rect 5448 9333 5457 9367
rect 5457 9333 5491 9367
rect 5491 9333 5500 9367
rect 5448 9324 5500 9333
rect 7380 9392 7432 9444
rect 7564 9392 7616 9444
rect 7012 9367 7064 9376
rect 7012 9333 7021 9367
rect 7021 9333 7055 9367
rect 7055 9333 7064 9367
rect 7012 9324 7064 9333
rect 7104 9367 7156 9376
rect 7104 9333 7113 9367
rect 7113 9333 7147 9367
rect 7147 9333 7156 9367
rect 7104 9324 7156 9333
rect 7748 9324 7800 9376
rect 9680 9324 9732 9376
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 6368 9120 6420 9172
rect 7472 9120 7524 9172
rect 10324 9120 10376 9172
rect 2044 9052 2096 9104
rect 3516 9052 3568 9104
rect 5448 9052 5500 9104
rect 4252 9027 4304 9036
rect 4252 8993 4261 9027
rect 4261 8993 4295 9027
rect 4295 8993 4304 9027
rect 4252 8984 4304 8993
rect 6828 9052 6880 9104
rect 7104 8984 7156 9036
rect 7380 9052 7432 9104
rect 9128 8984 9180 9036
rect 3608 8959 3660 8968
rect 3608 8925 3617 8959
rect 3617 8925 3651 8959
rect 3651 8925 3660 8959
rect 3608 8916 3660 8925
rect 9772 8916 9824 8968
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 2780 8780 2832 8832
rect 4896 8780 4948 8832
rect 7104 8780 7156 8832
rect 8668 8823 8720 8832
rect 8668 8789 8677 8823
rect 8677 8789 8711 8823
rect 8711 8789 8720 8823
rect 8668 8780 8720 8789
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 1768 8576 1820 8628
rect 4160 8576 4212 8628
rect 7564 8576 7616 8628
rect 9772 8619 9824 8628
rect 9772 8585 9781 8619
rect 9781 8585 9815 8619
rect 9815 8585 9824 8619
rect 9772 8576 9824 8585
rect 6276 8508 6328 8560
rect 4252 8440 4304 8492
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 388 8372 440 8424
rect 1216 8372 1268 8424
rect 1492 8372 1544 8424
rect 2688 8372 2740 8424
rect 4896 8372 4948 8424
rect 6552 8415 6604 8424
rect 6552 8381 6561 8415
rect 6561 8381 6595 8415
rect 6595 8381 6604 8415
rect 6552 8372 6604 8381
rect 8392 8415 8444 8424
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 3056 8304 3108 8356
rect 7104 8347 7156 8356
rect 7104 8313 7138 8347
rect 7138 8313 7156 8347
rect 7104 8304 7156 8313
rect 8116 8304 8168 8356
rect 1124 8236 1176 8288
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 2964 8236 3016 8245
rect 8208 8279 8260 8288
rect 8208 8245 8217 8279
rect 8217 8245 8251 8279
rect 8251 8245 8260 8279
rect 8208 8236 8260 8245
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 2688 8075 2740 8084
rect 2688 8041 2697 8075
rect 2697 8041 2731 8075
rect 2731 8041 2740 8075
rect 2688 8032 2740 8041
rect 7012 8032 7064 8084
rect 8392 8032 8444 8084
rect 8760 8032 8812 8084
rect 7104 7896 7156 7948
rect 6000 7692 6052 7744
rect 7288 7692 7340 7744
rect 8668 7896 8720 7948
rect 9220 7735 9272 7744
rect 9220 7701 9229 7735
rect 9229 7701 9263 7735
rect 9263 7701 9272 7735
rect 9220 7692 9272 7701
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 7104 7488 7156 7540
rect 2688 7352 2740 7404
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 1124 7327 1176 7336
rect 1124 7293 1158 7327
rect 1158 7293 1176 7327
rect 1124 7284 1176 7293
rect 3332 7284 3384 7336
rect 6000 7327 6052 7336
rect 6000 7293 6009 7327
rect 6009 7293 6043 7327
rect 6043 7293 6052 7327
rect 6000 7284 6052 7293
rect 7748 7284 7800 7336
rect 7840 7216 7892 7268
rect 8760 7284 8812 7336
rect 9496 7216 9548 7268
rect 2136 7148 2188 7200
rect 2872 7148 2924 7200
rect 4712 7191 4764 7200
rect 4712 7157 4721 7191
rect 4721 7157 4755 7191
rect 4755 7157 4764 7191
rect 4712 7148 4764 7157
rect 6000 7148 6052 7200
rect 6552 7148 6604 7200
rect 8484 7191 8536 7200
rect 8484 7157 8493 7191
rect 8493 7157 8527 7191
rect 8527 7157 8536 7191
rect 8484 7148 8536 7157
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 9220 6876 9272 6928
rect 2780 6808 2832 6860
rect 2872 6851 2924 6860
rect 2872 6817 2881 6851
rect 2881 6817 2915 6851
rect 2915 6817 2924 6851
rect 2872 6808 2924 6817
rect 4712 6808 4764 6860
rect 8760 6851 8812 6860
rect 8760 6817 8769 6851
rect 8769 6817 8803 6851
rect 8803 6817 8812 6851
rect 8760 6808 8812 6817
rect 9864 6851 9916 6860
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 2688 6740 2740 6792
rect 1860 6604 1912 6656
rect 9588 6672 9640 6724
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 4988 6647 5040 6656
rect 4988 6613 4997 6647
rect 4997 6613 5031 6647
rect 5031 6613 5040 6647
rect 4988 6604 5040 6613
rect 7748 6604 7800 6656
rect 8852 6647 8904 6656
rect 8852 6613 8861 6647
rect 8861 6613 8895 6647
rect 8895 6613 8904 6647
rect 8852 6604 8904 6613
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 7196 6400 7248 6452
rect 3976 6332 4028 6384
rect 6920 6332 6972 6384
rect 7380 6332 7432 6384
rect 2228 6196 2280 6248
rect 2964 6196 3016 6248
rect 6092 6239 6144 6248
rect 6092 6205 6101 6239
rect 6101 6205 6135 6239
rect 6135 6205 6144 6239
rect 6092 6196 6144 6205
rect 6368 6239 6420 6248
rect 6368 6205 6377 6239
rect 6377 6205 6411 6239
rect 6411 6205 6420 6239
rect 6368 6196 6420 6205
rect 6552 6239 6604 6248
rect 6552 6205 6561 6239
rect 6561 6205 6595 6239
rect 6595 6205 6604 6239
rect 6552 6196 6604 6205
rect 3240 6060 3292 6112
rect 5816 6171 5868 6180
rect 5816 6137 5825 6171
rect 5825 6137 5859 6171
rect 5859 6137 5868 6171
rect 5816 6128 5868 6137
rect 6184 6060 6236 6112
rect 7196 6128 7248 6180
rect 7472 6239 7524 6248
rect 7472 6205 7481 6239
rect 7481 6205 7515 6239
rect 7515 6205 7524 6239
rect 7472 6196 7524 6205
rect 8760 6400 8812 6452
rect 9864 6400 9916 6452
rect 7656 6128 7708 6180
rect 7564 6103 7616 6112
rect 7564 6069 7573 6103
rect 7573 6069 7607 6103
rect 7607 6069 7616 6103
rect 7564 6060 7616 6069
rect 8852 6060 8904 6112
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 5816 5856 5868 5908
rect 7656 5856 7708 5908
rect 9128 5899 9180 5908
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 9496 5856 9548 5908
rect 2320 5788 2372 5840
rect 3332 5788 3384 5840
rect 3976 5788 4028 5840
rect 4160 5720 4212 5772
rect 7472 5788 7524 5840
rect 1768 5652 1820 5704
rect 4252 5695 4304 5704
rect 4252 5661 4261 5695
rect 4261 5661 4295 5695
rect 4295 5661 4304 5695
rect 4252 5652 4304 5661
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 6092 5720 6144 5772
rect 5632 5584 5684 5636
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 7196 5763 7248 5772
rect 7196 5729 7205 5763
rect 7205 5729 7239 5763
rect 7239 5729 7248 5763
rect 7196 5720 7248 5729
rect 7380 5720 7432 5772
rect 7564 5652 7616 5704
rect 9680 5720 9732 5772
rect 6828 5584 6880 5636
rect 7012 5516 7064 5568
rect 8392 5516 8444 5568
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 8392 5355 8444 5364
rect 8392 5321 8401 5355
rect 8401 5321 8435 5355
rect 8435 5321 8444 5355
rect 8392 5312 8444 5321
rect 3148 5108 3200 5160
rect 3332 5176 3384 5228
rect 5540 5176 5592 5228
rect 7288 5176 7340 5228
rect 9128 5176 9180 5228
rect 3424 5151 3476 5160
rect 3424 5117 3433 5151
rect 3433 5117 3467 5151
rect 3467 5117 3476 5151
rect 3424 5108 3476 5117
rect 5632 5108 5684 5160
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 2688 5083 2740 5092
rect 2688 5049 2697 5083
rect 2697 5049 2731 5083
rect 2731 5049 2740 5083
rect 2688 5040 2740 5049
rect 2964 5040 3016 5092
rect 5356 5040 5408 5092
rect 7012 5083 7064 5092
rect 7012 5049 7021 5083
rect 7021 5049 7055 5083
rect 7055 5049 7064 5083
rect 7012 5040 7064 5049
rect 2320 4972 2372 5024
rect 4712 4972 4764 5024
rect 6092 4972 6144 5024
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 4160 4811 4212 4820
rect 4160 4777 4169 4811
rect 4169 4777 4203 4811
rect 4203 4777 4212 4811
rect 4160 4768 4212 4777
rect 1768 4700 1820 4752
rect 2780 4700 2832 4752
rect 3148 4700 3200 4752
rect 3332 4700 3384 4752
rect 4068 4700 4120 4752
rect 1216 4675 1268 4684
rect 1216 4641 1250 4675
rect 1250 4641 1268 4675
rect 1216 4632 1268 4641
rect 3240 4675 3292 4684
rect 3240 4641 3249 4675
rect 3249 4641 3283 4675
rect 3283 4641 3292 4675
rect 3240 4632 3292 4641
rect 4712 4768 4764 4820
rect 4804 4768 4856 4820
rect 5632 4768 5684 4820
rect 6920 4811 6972 4820
rect 6920 4777 6929 4811
rect 6929 4777 6963 4811
rect 6963 4777 6972 4811
rect 6920 4768 6972 4777
rect 4528 4743 4580 4752
rect 4528 4709 4537 4743
rect 4537 4709 4571 4743
rect 4571 4709 4580 4743
rect 4528 4700 4580 4709
rect 4988 4700 5040 4752
rect 5724 4700 5776 4752
rect 3424 4564 3476 4616
rect 4804 4632 4856 4684
rect 4896 4564 4948 4616
rect 2872 4471 2924 4480
rect 2872 4437 2881 4471
rect 2881 4437 2915 4471
rect 2915 4437 2924 4471
rect 2872 4428 2924 4437
rect 5264 4428 5316 4480
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 6092 4675 6144 4684
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 6276 4632 6328 4684
rect 7656 4632 7708 4684
rect 7748 4675 7800 4684
rect 7748 4641 7757 4675
rect 7757 4641 7791 4675
rect 7791 4641 7800 4675
rect 7748 4632 7800 4641
rect 8484 4632 8536 4684
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 7472 4564 7524 4616
rect 8208 4564 8260 4616
rect 9772 4564 9824 4616
rect 7564 4496 7616 4548
rect 6828 4428 6880 4480
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 2872 4267 2924 4276
rect 2872 4233 2881 4267
rect 2881 4233 2915 4267
rect 2915 4233 2924 4267
rect 2872 4224 2924 4233
rect 5816 4224 5868 4276
rect 5632 4156 5684 4208
rect 4252 4088 4304 4140
rect 4988 4088 5040 4140
rect 1768 4020 1820 4072
rect 2136 3952 2188 4004
rect 1216 3884 1268 3936
rect 2596 3927 2648 3936
rect 2596 3893 2605 3927
rect 2605 3893 2639 3927
rect 2639 3893 2648 3927
rect 2596 3884 2648 3893
rect 2964 3952 3016 4004
rect 3240 4063 3292 4072
rect 3240 4029 3249 4063
rect 3249 4029 3283 4063
rect 3283 4029 3292 4063
rect 3240 4020 3292 4029
rect 4068 4020 4120 4072
rect 5540 4020 5592 4072
rect 5724 4020 5776 4072
rect 3884 3884 3936 3936
rect 4160 3952 4212 4004
rect 4804 3952 4856 4004
rect 6092 4063 6144 4072
rect 6092 4029 6101 4063
rect 6101 4029 6135 4063
rect 6135 4029 6144 4063
rect 6092 4020 6144 4029
rect 8024 4088 8076 4140
rect 6276 4020 6328 4072
rect 6460 4063 6512 4072
rect 6460 4029 6469 4063
rect 6469 4029 6503 4063
rect 6503 4029 6512 4063
rect 6460 4020 6512 4029
rect 6552 4020 6604 4072
rect 7196 4063 7248 4072
rect 7196 4029 7205 4063
rect 7205 4029 7239 4063
rect 7239 4029 7248 4063
rect 7196 4020 7248 4029
rect 7380 4020 7432 4072
rect 7472 4063 7524 4072
rect 7472 4029 7481 4063
rect 7481 4029 7515 4063
rect 7515 4029 7524 4063
rect 7472 4020 7524 4029
rect 7656 4020 7708 4072
rect 8116 4020 8168 4072
rect 4252 3884 4304 3936
rect 6276 3884 6328 3936
rect 7564 3884 7616 3936
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 2964 3680 3016 3732
rect 3332 3680 3384 3732
rect 3424 3723 3476 3732
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 4896 3680 4948 3732
rect 6184 3680 6236 3732
rect 7196 3680 7248 3732
rect 7288 3680 7340 3732
rect 8300 3680 8352 3732
rect 8760 3680 8812 3732
rect 2044 3587 2096 3596
rect 2044 3553 2053 3587
rect 2053 3553 2087 3587
rect 2087 3553 2096 3587
rect 2044 3544 2096 3553
rect 2596 3544 2648 3596
rect 3056 3544 3108 3596
rect 3240 3544 3292 3596
rect 3976 3655 4028 3664
rect 3976 3621 3985 3655
rect 3985 3621 4019 3655
rect 4019 3621 4028 3655
rect 3976 3612 4028 3621
rect 4160 3612 4212 3664
rect 5632 3612 5684 3664
rect 2136 3451 2188 3460
rect 2136 3417 2145 3451
rect 2145 3417 2179 3451
rect 2179 3417 2188 3451
rect 2136 3408 2188 3417
rect 2320 3383 2372 3392
rect 2320 3349 2329 3383
rect 2329 3349 2363 3383
rect 2363 3349 2372 3383
rect 2320 3340 2372 3349
rect 2780 3519 2832 3528
rect 2780 3485 2789 3519
rect 2789 3485 2823 3519
rect 2823 3485 2832 3519
rect 2780 3476 2832 3485
rect 3424 3476 3476 3528
rect 3516 3476 3568 3528
rect 6460 3544 6512 3596
rect 7012 3544 7064 3596
rect 7104 3587 7156 3596
rect 7104 3553 7113 3587
rect 7113 3553 7147 3587
rect 7147 3553 7156 3587
rect 7104 3544 7156 3553
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 4252 3476 4304 3485
rect 7288 3587 7340 3596
rect 7288 3553 7297 3587
rect 7297 3553 7331 3587
rect 7331 3553 7340 3587
rect 7288 3544 7340 3553
rect 8392 3476 8444 3528
rect 3056 3408 3108 3460
rect 3240 3451 3292 3460
rect 3240 3417 3249 3451
rect 3249 3417 3283 3451
rect 3283 3417 3292 3451
rect 3240 3408 3292 3417
rect 5264 3408 5316 3460
rect 6092 3408 6144 3460
rect 2780 3340 2832 3392
rect 8484 3340 8536 3392
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 3516 3136 3568 3188
rect 4712 3136 4764 3188
rect 5080 3136 5132 3188
rect 7104 3136 7156 3188
rect 7748 3136 7800 3188
rect 8024 3179 8076 3188
rect 8024 3145 8033 3179
rect 8033 3145 8067 3179
rect 8067 3145 8076 3179
rect 8024 3136 8076 3145
rect 9496 3136 9548 3188
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 4804 3111 4856 3120
rect 4804 3077 4813 3111
rect 4813 3077 4847 3111
rect 4847 3077 4856 3111
rect 4804 3068 4856 3077
rect 7380 3068 7432 3120
rect 7288 3000 7340 3052
rect 4252 2932 4304 2984
rect 4896 2932 4948 2984
rect 5172 2932 5224 2984
rect 3516 2907 3568 2916
rect 3516 2873 3550 2907
rect 3550 2873 3568 2907
rect 3516 2864 3568 2873
rect 4988 2864 5040 2916
rect 5264 2907 5316 2916
rect 5264 2873 5273 2907
rect 5273 2873 5307 2907
rect 5307 2873 5316 2907
rect 5264 2864 5316 2873
rect 8300 3000 8352 3052
rect 5632 2839 5684 2848
rect 5632 2805 5641 2839
rect 5641 2805 5675 2839
rect 5675 2805 5684 2839
rect 5632 2796 5684 2805
rect 8024 2839 8076 2848
rect 8024 2805 8051 2839
rect 8051 2805 8076 2839
rect 8024 2796 8076 2805
rect 8208 2907 8260 2916
rect 8208 2873 8217 2907
rect 8217 2873 8251 2907
rect 8251 2873 8260 2907
rect 8208 2864 8260 2873
rect 8484 2932 8536 2984
rect 8760 2864 8812 2916
rect 8392 2796 8444 2848
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 4988 2592 5040 2644
rect 3148 2524 3200 2576
rect 2780 2456 2832 2508
rect 4068 2524 4120 2576
rect 6092 2592 6144 2644
rect 6368 2592 6420 2644
rect 7012 2592 7064 2644
rect 5172 2456 5224 2508
rect 5264 2388 5316 2440
rect 5632 2499 5684 2508
rect 5632 2465 5641 2499
rect 5641 2465 5675 2499
rect 5675 2465 5684 2499
rect 5632 2456 5684 2465
rect 7840 2524 7892 2576
rect 7932 2567 7984 2576
rect 7932 2533 7941 2567
rect 7941 2533 7975 2567
rect 7975 2533 7984 2567
rect 7932 2524 7984 2533
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 7748 2499 7800 2508
rect 7748 2465 7757 2499
rect 7757 2465 7791 2499
rect 7791 2465 7800 2499
rect 7748 2456 7800 2465
rect 8024 2499 8076 2508
rect 8024 2465 8033 2499
rect 8033 2465 8067 2499
rect 8067 2465 8076 2499
rect 8024 2456 8076 2465
rect 8208 2456 8260 2508
rect 4804 2320 4856 2372
rect 4712 2252 4764 2304
rect 5540 2295 5592 2304
rect 5540 2261 5549 2295
rect 5549 2261 5583 2295
rect 5583 2261 5592 2295
rect 5540 2252 5592 2261
rect 7012 2252 7064 2304
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 5264 2048 5316 2100
rect 7840 2048 7892 2100
rect 8760 2091 8812 2100
rect 8760 2057 8769 2091
rect 8769 2057 8803 2091
rect 8803 2057 8812 2091
rect 8760 2048 8812 2057
rect 4252 1955 4304 1964
rect 4252 1921 4261 1955
rect 4261 1921 4295 1955
rect 4295 1921 4304 1955
rect 4252 1912 4304 1921
rect 5632 1844 5684 1896
rect 6092 1887 6144 1896
rect 6092 1853 6101 1887
rect 6101 1853 6135 1887
rect 6135 1853 6144 1887
rect 6092 1844 6144 1853
rect 4252 1776 4304 1828
rect 6920 1980 6972 2032
rect 7012 1912 7064 1964
rect 6920 1887 6972 1896
rect 6920 1853 6929 1887
rect 6929 1853 6963 1887
rect 6963 1853 6972 1887
rect 6920 1844 6972 1853
rect 7932 1912 7984 1964
rect 7932 1776 7984 1828
rect 8024 1819 8076 1828
rect 8024 1785 8033 1819
rect 8033 1785 8067 1819
rect 8067 1785 8076 1819
rect 8024 1776 8076 1785
rect 8392 1887 8444 1896
rect 8392 1853 8401 1887
rect 8401 1853 8435 1887
rect 8435 1853 8444 1887
rect 8392 1844 8444 1853
rect 9772 1912 9824 1964
rect 6736 1751 6788 1760
rect 6736 1717 6745 1751
rect 6745 1717 6779 1751
rect 6779 1717 6788 1751
rect 6736 1708 6788 1717
rect 7564 1751 7616 1760
rect 7564 1717 7573 1751
rect 7573 1717 7607 1751
rect 7607 1717 7616 1751
rect 7564 1708 7616 1717
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 4252 1504 4304 1556
rect 4712 1547 4764 1556
rect 4712 1513 4739 1547
rect 4739 1513 4764 1547
rect 4712 1504 4764 1513
rect 6092 1504 6144 1556
rect 4068 1436 4120 1488
rect 6828 1504 6880 1556
rect 7932 1504 7984 1556
rect 6736 1436 6788 1488
rect 8300 1436 8352 1488
rect 7564 1411 7616 1420
rect 7564 1377 7598 1411
rect 7598 1377 7616 1411
rect 7564 1368 7616 1377
rect 5540 1164 5592 1216
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
<< metal2 >>
rect 386 9957 442 10757
rect 1214 9957 1270 10757
rect 2042 9957 2098 10757
rect 2870 9957 2926 10757
rect 3698 9957 3754 10757
rect 4526 9957 4582 10757
rect 5354 9957 5410 10757
rect 6182 9957 6238 10757
rect 7010 9957 7066 10757
rect 7838 9957 7894 10757
rect 8666 9957 8722 10757
rect 9494 9957 9550 10757
rect 10322 9957 10378 10757
rect 400 8430 428 9957
rect 1228 8430 1256 9957
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 9178 1624 9454
rect 1768 9444 1820 9450
rect 1768 9386 1820 9392
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1504 8430 1532 8774
rect 1780 8634 1808 9386
rect 2056 9110 2084 9957
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 2700 8430 2728 9522
rect 2884 9518 2912 9957
rect 3712 9926 3740 9957
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3528 9518 3556 9862
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 4540 9722 4568 9957
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 5368 9518 5396 9957
rect 6196 9654 6224 9957
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 388 8424 440 8430
rect 388 8366 440 8372
rect 1216 8424 1268 8430
rect 1216 8366 1268 8372
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 1124 8288 1176 8294
rect 1124 8230 1176 8236
rect 1136 7342 1164 8230
rect 2700 8090 2728 8366
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2700 7410 2728 8026
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 1124 7336 1176 7342
rect 1124 7278 1176 7284
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2148 6914 2176 7142
rect 2148 6886 2268 6914
rect 2240 6798 2268 6886
rect 2700 6798 2728 7346
rect 2792 6866 2820 8774
rect 3068 8362 3096 9318
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2884 6866 2912 7142
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1768 5704 1820 5710
rect 1872 5692 1900 6598
rect 2240 6254 2268 6734
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2332 5846 2360 6598
rect 2976 6254 3004 8230
rect 3344 7342 3372 9318
rect 3528 9110 3556 9318
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3620 8974 3648 9318
rect 4264 9042 4292 9386
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 4322 9276 4630 9285
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 5460 9110 5488 9318
rect 6380 9178 6408 9454
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 1820 5664 1900 5692
rect 1768 5646 1820 5652
rect 1780 4758 1808 5646
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 2688 5092 2740 5098
rect 2688 5034 2740 5040
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 1768 4752 1820 4758
rect 1768 4694 1820 4700
rect 1216 4684 1268 4690
rect 1216 4626 1268 4632
rect 1228 3942 1256 4626
rect 1780 4078 1808 4694
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 2136 4004 2188 4010
rect 2136 3946 2188 3952
rect 1216 3936 1268 3942
rect 1216 3878 1268 3884
rect 2042 3632 2098 3641
rect 2042 3567 2044 3576
rect 2096 3567 2098 3576
rect 2044 3538 2096 3544
rect 2148 3466 2176 3946
rect 2136 3460 2188 3466
rect 2136 3402 2188 3408
rect 2332 3398 2360 4966
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2608 3602 2636 3878
rect 2700 3641 2728 5034
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 2686 3632 2742 3641
rect 2596 3596 2648 3602
rect 2686 3567 2742 3576
rect 2596 3538 2648 3544
rect 2792 3534 2820 4694
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2884 4282 2912 4422
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2976 4010 3004 5034
rect 3160 4758 3188 5102
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2976 3738 3004 3946
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 3068 3466 3096 3538
rect 3160 3482 3188 4694
rect 3252 4690 3280 6054
rect 3988 5846 4016 6326
rect 4172 5930 4200 8570
rect 4264 8498 4292 8978
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4908 8430 4936 8774
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6012 7342 6040 7686
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 4724 6866 4752 7142
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 4080 5902 4200 5930
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 3344 5234 3372 5782
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3332 4752 3384 4758
rect 3332 4694 3384 4700
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3344 4570 3372 4694
rect 3436 4622 3464 5102
rect 4080 4758 4108 5902
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4172 4826 4200 5714
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 3252 4542 3372 4570
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3252 4078 3280 4542
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3252 3602 3280 4014
rect 3436 3738 3464 4558
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 4080 4078 4108 4694
rect 4264 4146 4292 5646
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 4724 4826 4752 4966
rect 4816 4826 4844 5646
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4528 4752 4580 4758
rect 4526 4720 4528 4729
rect 4580 4720 4582 4729
rect 4526 4655 4582 4664
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 3884 3936 3936 3942
rect 3936 3896 4108 3924
rect 3884 3878 3936 3884
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3160 3466 3280 3482
rect 3056 3460 3108 3466
rect 3160 3460 3292 3466
rect 3160 3454 3240 3460
rect 3056 3402 3108 3408
rect 3240 3402 3292 3408
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2792 2514 2820 3334
rect 3344 2774 3372 3674
rect 3436 3534 3464 3674
rect 3976 3664 4028 3670
rect 3974 3632 3976 3641
rect 4028 3632 4030 3641
rect 3974 3567 4030 3576
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3528 3194 3556 3470
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3160 2746 3372 2774
rect 3160 2582 3188 2746
rect 3528 2650 3556 2858
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 4080 2582 4108 3896
rect 4172 3670 4200 3946
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 4264 3534 4292 3878
rect 4322 3836 4630 3845
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4264 2990 4292 3470
rect 4724 3194 4752 4762
rect 5000 4758 5028 6598
rect 5816 6180 5868 6186
rect 5816 6122 5868 6128
rect 5828 5914 5856 6122
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 4988 4752 5040 4758
rect 4988 4694 5040 4700
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4816 4010 4844 4626
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 4908 3738 4936 4558
rect 5000 4146 5028 4694
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 4068 2576 4120 2582
rect 4068 2518 4120 2524
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 4080 1494 4108 2518
rect 4264 1970 4292 2926
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 4816 2378 4844 3062
rect 4908 2990 4936 3674
rect 5276 3466 5304 4422
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 5000 2650 5028 2858
rect 5092 2825 5120 3130
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5078 2816 5134 2825
rect 5078 2751 5134 2760
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5184 2514 5212 2926
rect 5276 2922 5304 3402
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 5262 2816 5318 2825
rect 5262 2751 5318 2760
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 5276 2446 5304 2751
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 4804 2372 4856 2378
rect 4804 2314 4856 2320
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 4252 1964 4304 1970
rect 4252 1906 4304 1912
rect 4252 1828 4304 1834
rect 4252 1770 4304 1776
rect 4264 1562 4292 1770
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 4724 1562 4752 2246
rect 5276 2106 5304 2382
rect 5264 2100 5316 2106
rect 5264 2042 5316 2048
rect 4252 1556 4304 1562
rect 4252 1498 4304 1504
rect 4712 1556 4764 1562
rect 4712 1498 4764 1504
rect 4068 1488 4120 1494
rect 4068 1430 4120 1436
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 5368 800 5396 5034
rect 5552 4078 5580 5170
rect 5644 5166 5672 5578
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5644 4826 5672 5102
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5724 4752 5776 4758
rect 6012 4729 6040 7142
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6104 5778 6132 6190
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6196 5710 6224 6054
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 5724 4694 5776 4700
rect 5998 4720 6054 4729
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5644 3670 5672 4150
rect 5736 4078 5764 4694
rect 5816 4684 5868 4690
rect 6104 4690 6132 4966
rect 6288 4690 6316 8502
rect 6564 8430 6592 9658
rect 7024 9586 7052 9957
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6840 8498 6868 9046
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6840 7970 6868 8434
rect 7024 8090 7052 9318
rect 7116 9042 7144 9318
rect 7392 9110 7420 9386
rect 7484 9178 7512 9454
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 8362 7144 8774
rect 7576 8634 7604 9386
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 6840 7954 7144 7970
rect 6840 7948 7156 7954
rect 6840 7942 7104 7948
rect 7104 7890 7156 7896
rect 7116 7546 7144 7890
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 6254 6592 7142
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 5998 4655 6000 4664
rect 5816 4626 5868 4632
rect 6052 4655 6054 4664
rect 6092 4684 6144 4690
rect 6000 4626 6052 4632
rect 6092 4626 6144 4632
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 5828 4282 5856 4626
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5724 4072 5776 4078
rect 6092 4072 6144 4078
rect 5724 4014 5776 4020
rect 6090 4040 6092 4049
rect 6144 4040 6146 4049
rect 6090 3975 6146 3984
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 6104 3466 6132 3975
rect 6196 3738 6224 4558
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6288 3942 6316 4014
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5644 2514 5672 2790
rect 6380 2650 6408 6190
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6840 5166 6868 5578
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6840 4486 6868 5102
rect 6932 4826 6960 6326
rect 7208 6186 7236 6394
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7024 5574 7052 5646
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7012 5092 7064 5098
rect 7208 5080 7236 5714
rect 7300 5234 7328 7686
rect 7760 7342 7788 9318
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7852 7274 7880 9957
rect 8680 9722 8708 9957
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8404 8430 8432 9454
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8128 7546 8156 8298
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7392 5778 7420 6326
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7484 5846 7512 6190
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7576 5710 7604 6054
rect 7668 5914 7696 6122
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7064 5052 7236 5080
rect 7012 5034 7064 5040
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6460 4072 6512 4078
rect 6552 4072 6604 4078
rect 6460 4014 6512 4020
rect 6550 4040 6552 4049
rect 6604 4040 6606 4049
rect 6472 3602 6500 4014
rect 6550 3975 6606 3984
rect 7024 3602 7052 5034
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7208 3738 7236 4014
rect 7300 3738 7328 5170
rect 7760 4690 7788 6598
rect 8220 4706 8248 8230
rect 8404 8090 8432 8366
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8680 7954 8708 8774
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8772 7342 8800 8026
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8404 5370 8432 5510
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 8128 4678 8248 4706
rect 8496 4690 8524 7142
rect 8772 6866 8800 7278
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8484 4684 8536 4690
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7484 4078 7512 4558
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7024 2650 7052 3538
rect 7116 3194 7144 3538
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7300 3058 7328 3538
rect 7392 3126 7420 4014
rect 7576 3942 7604 4490
rect 7668 4078 7696 4626
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 8036 3194 8064 4082
rect 8128 4078 8156 4678
rect 8484 4626 8536 4632
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5552 1222 5580 2246
rect 5644 1902 5672 2450
rect 6104 1902 6132 2586
rect 7024 2394 7052 2586
rect 7760 2514 7788 3130
rect 8220 2938 8248 4558
rect 8772 3738 8800 6394
rect 8864 6118 8892 6598
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 9140 5914 9168 8978
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9232 6934 9260 7686
rect 9508 7392 9536 9957
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9508 7364 9628 7392
rect 9496 7268 9548 7274
rect 9496 7210 9548 7216
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 9508 5914 9536 7210
rect 9600 6730 9628 7364
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9140 5234 9168 5850
rect 9692 5778 9720 9318
rect 10336 9178 10364 9957
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9784 8634 9812 8910
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9876 6458 9904 6802
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8312 3058 8340 3674
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 7944 2922 8248 2938
rect 7944 2916 8260 2922
rect 7944 2910 8208 2916
rect 7944 2582 7972 2910
rect 8208 2858 8260 2864
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 6932 2366 7052 2394
rect 6932 2038 6960 2366
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 6920 2032 6972 2038
rect 6920 1974 6972 1980
rect 6932 1902 6960 1974
rect 7024 1970 7052 2246
rect 7852 2106 7880 2518
rect 7840 2100 7892 2106
rect 7840 2042 7892 2048
rect 7944 1970 7972 2518
rect 8036 2514 8064 2790
rect 8312 2530 8340 2994
rect 8404 2854 8432 3470
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8496 2990 8524 3334
rect 9784 3194 9812 4558
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8220 2514 8340 2530
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 8208 2508 8340 2514
rect 8260 2502 8340 2508
rect 8208 2450 8260 2456
rect 7012 1964 7064 1970
rect 7012 1906 7064 1912
rect 7932 1964 7984 1970
rect 7932 1906 7984 1912
rect 5632 1896 5684 1902
rect 5632 1838 5684 1844
rect 6092 1896 6144 1902
rect 6092 1838 6144 1844
rect 6920 1896 6972 1902
rect 6920 1838 6972 1844
rect 6104 1562 6132 1838
rect 6736 1760 6788 1766
rect 6736 1702 6788 1708
rect 6092 1556 6144 1562
rect 6092 1498 6144 1504
rect 6748 1494 6776 1702
rect 6932 1578 6960 1838
rect 7944 1834 7972 1906
rect 8036 1834 8064 2450
rect 7932 1828 7984 1834
rect 7932 1770 7984 1776
rect 8024 1828 8076 1834
rect 8024 1770 8076 1776
rect 7564 1760 7616 1766
rect 7564 1702 7616 1708
rect 6840 1562 6960 1578
rect 6828 1556 6960 1562
rect 6880 1550 6960 1556
rect 6828 1498 6880 1504
rect 6736 1488 6788 1494
rect 6736 1430 6788 1436
rect 7576 1426 7604 1702
rect 7944 1562 7972 1770
rect 7932 1556 7984 1562
rect 7932 1498 7984 1504
rect 8312 1494 8340 2502
rect 8404 1902 8432 2790
rect 8772 2106 8800 2858
rect 9508 2650 9536 3130
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 8760 2100 8812 2106
rect 8760 2042 8812 2048
rect 9784 1970 9812 3130
rect 9772 1964 9824 1970
rect 9772 1906 9824 1912
rect 8392 1896 8444 1902
rect 8392 1838 8444 1844
rect 8300 1488 8352 1494
rect 8300 1430 8352 1436
rect 7564 1420 7616 1426
rect 7564 1362 7616 1368
rect 5540 1216 5592 1222
rect 5540 1158 5592 1164
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
rect 5354 0 5410 800
<< via2 >>
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 2042 3596 2098 3632
rect 2042 3576 2044 3596
rect 2044 3576 2096 3596
rect 2096 3576 2098 3596
rect 2686 3576 2742 3632
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 4526 4700 4528 4720
rect 4528 4700 4580 4720
rect 4580 4700 4582 4720
rect 4526 4664 4582 4700
rect 3974 3612 3976 3632
rect 3976 3612 4028 3632
rect 4028 3612 4030 3632
rect 3974 3576 4030 3612
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 5078 2760 5134 2816
rect 5262 2760 5318 2816
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 5998 4684 6054 4720
rect 5998 4664 6000 4684
rect 6000 4664 6052 4684
rect 6052 4664 6054 4684
rect 6090 4020 6092 4040
rect 6092 4020 6144 4040
rect 6144 4020 6146 4040
rect 6090 3984 6146 4020
rect 6550 4020 6552 4040
rect 6552 4020 6604 4040
rect 6604 4020 6606 4040
rect 6550 3984 6606 4020
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
<< metal3 >>
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 4521 4722 4587 4725
rect 5993 4722 6059 4725
rect 4521 4720 6059 4722
rect 4521 4664 4526 4720
rect 4582 4664 5998 4720
rect 6054 4664 6059 4720
rect 4521 4662 6059 4664
rect 4521 4659 4587 4662
rect 5993 4659 6059 4662
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 6085 4042 6151 4045
rect 6545 4042 6611 4045
rect 6085 4040 6611 4042
rect 6085 3984 6090 4040
rect 6146 3984 6550 4040
rect 6606 3984 6611 4040
rect 6085 3982 6611 3984
rect 6085 3979 6151 3982
rect 6545 3979 6611 3982
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 4318 3775 4634 3776
rect 2037 3634 2103 3637
rect 2681 3634 2747 3637
rect 3969 3634 4035 3637
rect 2037 3632 4035 3634
rect 2037 3576 2042 3632
rect 2098 3576 2686 3632
rect 2742 3576 3974 3632
rect 4030 3576 4035 3632
rect 2037 3574 4035 3576
rect 2037 3571 2103 3574
rect 2681 3571 2747 3574
rect 3969 3571 4035 3574
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 5073 2818 5139 2821
rect 5257 2818 5323 2821
rect 5073 2816 5323 2818
rect 5073 2760 5078 2816
rect 5134 2760 5262 2816
rect 5318 2760 5323 2816
rect 5073 2758 5323 2760
rect 5073 2755 5139 2758
rect 5257 2755 5323 2758
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
<< via3 >>
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
<< metal4 >>
rect 3656 9824 3976 9840
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 9280 4636 9840
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4316 8192 4636 9216
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
use sky130_fd_sc_hd__inv_2  _054_
timestamp 28801
transform 1 0 3864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _055_
timestamp 28801
transform 1 0 7728 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp 28801
transform -1 0 6072 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 28801
transform 1 0 5980 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 28801
transform 1 0 9476 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _059_
timestamp 28801
transform -1 0 9384 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _060_
timestamp 28801
transform 1 0 5796 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _061_
timestamp 28801
transform 1 0 6348 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _062_
timestamp 28801
transform 1 0 6624 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _063_
timestamp 28801
transform -1 0 8004 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _064_
timestamp 28801
transform 1 0 3220 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _065_
timestamp 28801
transform 1 0 7084 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _066_
timestamp 28801
transform -1 0 9384 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _067_
timestamp 28801
transform -1 0 6440 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _068_
timestamp 28801
transform -1 0 7268 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _069_
timestamp 28801
transform 1 0 3772 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _070_
timestamp 28801
transform 1 0 3220 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _071_
timestamp 28801
transform 1 0 3036 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _072_
timestamp 28801
transform 1 0 4232 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _073_
timestamp 28801
transform 1 0 4232 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _074_
timestamp 28801
transform 1 0 6624 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _075_
timestamp 28801
transform 1 0 5796 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _076_
timestamp 28801
transform -1 0 7728 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _077_
timestamp 28801
transform -1 0 6900 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _078_
timestamp 28801
transform -1 0 7820 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _079_
timestamp 28801
transform 1 0 5796 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _080_
timestamp 28801
transform 1 0 2484 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _081_
timestamp 28801
transform -1 0 3496 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _082_
timestamp 28801
transform -1 0 3128 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _083_
timestamp 28801
transform -1 0 2944 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _084_
timestamp 28801
transform 1 0 1840 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _085_
timestamp 28801
transform -1 0 2576 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _086_
timestamp 28801
transform 1 0 3220 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _087_
timestamp 28801
transform 1 0 4692 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _088_
timestamp 28801
transform -1 0 3220 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _089_
timestamp 28801
transform -1 0 3956 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _090_
timestamp 28801
transform -1 0 5704 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _091_
timestamp 28801
transform -1 0 7728 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _092_
timestamp 28801
transform 1 0 5244 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _093_
timestamp 28801
transform -1 0 5704 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _094_
timestamp 28801
transform 1 0 4876 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _095_
timestamp 28801
transform -1 0 4968 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _096_
timestamp 28801
transform 1 0 5888 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _097_
timestamp 28801
transform 1 0 5888 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _098_
timestamp 28801
transform -1 0 7084 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _099_
timestamp 28801
transform 1 0 6348 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _100_
timestamp 28801
transform -1 0 8096 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _101_
timestamp 28801
transform -1 0 7636 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _102_
timestamp 28801
transform 1 0 7544 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _103_
timestamp 28801
transform -1 0 8280 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 28801
transform 1 0 8372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _105_
timestamp 28801
transform 1 0 7084 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _106_
timestamp 28801
transform -1 0 7820 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _107_
timestamp 28801
transform -1 0 7636 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _108_
timestamp 28801
transform 1 0 7728 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _109_
timestamp 28801
transform 1 0 8372 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _110_
timestamp 28801
transform -1 0 5796 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _111_
timestamp 28801
transform 1 0 920 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _112_
timestamp 28801
transform 1 0 1196 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _113_
timestamp 28801
transform 1 0 3220 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _114_
timestamp 28801
transform 1 0 4232 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _115_
timestamp 28801
transform 1 0 4232 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _116_
timestamp 28801
transform -1 0 7268 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _117_
timestamp 28801
transform 1 0 7268 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _118_
timestamp 28801
transform 1 0 8096 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _119_
timestamp 28801
transform 1 0 8372 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _120_
timestamp 28801
transform 1 0 828 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _121_
timestamp 28801
transform 1 0 1840 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _122_
timestamp 28801
transform -1 0 2300 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _123_
timestamp 28801
transform -1 0 2300 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _124_
timestamp 28801
transform 1 0 3220 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _125_
timestamp 28801
transform -1 0 3036 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _126_
timestamp 28801
transform -1 0 5244 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _127_
timestamp 28801
transform 1 0 4232 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _128_
timestamp 28801
transform 1 0 5796 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _129_
timestamp 28801
transform 1 0 7268 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _130_
timestamp 28801
transform 1 0 8372 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _131_
timestamp 28801
transform 1 0 8372 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _132_
timestamp 28801
transform 1 0 1564 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _133_
timestamp 28801
transform 1 0 1656 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _134_
timestamp 28801
transform 1 0 3588 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _135_
timestamp 28801
transform 1 0 3220 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _136_
timestamp 28801
transform 1 0 4784 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _137_
timestamp 28801
transform -1 0 7268 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _138_
timestamp 28801
transform -1 0 7912 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _139_
timestamp 28801
transform -1 0 8832 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _140_
timestamp 28801
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _141_
timestamp 28801
transform -1 0 9936 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK
timestamp 28801
transform 1 0 4784 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_CLK
timestamp 28801
transform -1 0 5336 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_CLK
timestamp 28801
transform 1 0 7636 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_CLK
timestamp 28801
transform -1 0 4048 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_CLK
timestamp 28801
transform 1 0 7360 0 -1 8160
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636997256
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636997256
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 28801
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636997256
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636997256
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 28801
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636997256
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636997256
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 28801
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636997256
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_97
timestamp 28801
transform 1 0 9476 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_101
timestamp 28801
transform 1 0 9844 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636997256
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636997256
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636997256
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_39
timestamp 28801
transform 1 0 4140 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_48
timestamp 28801
transform 1 0 4968 0 -1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_89
timestamp 1636997256
transform 1 0 8740 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_101
timestamp 28801
transform 1 0 9844 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636997256
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636997256
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 28801
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 28801
transform 1 0 3220 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_37
timestamp 28801
transform 1 0 3956 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_56
timestamp 28801
transform 1 0 5704 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_68
timestamp 28801
transform 1 0 6808 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 28801
transform 1 0 8096 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_88
timestamp 28801
transform 1 0 8648 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_100
timestamp 28801
transform 1 0 9752 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636997256
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636997256
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_27
timestamp 28801
transform 1 0 3036 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_31
timestamp 28801
transform 1 0 3404 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_37
timestamp 28801
transform 1 0 3956 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_45
timestamp 28801
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 28801
transform 1 0 5796 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_65
timestamp 28801
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_98
timestamp 28801
transform 1 0 9568 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636997256
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636997256
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 28801
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_48
timestamp 28801
transform 1 0 4968 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_56
timestamp 1636997256
transform 1 0 5704 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_68
timestamp 28801
transform 1 0 6808 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_101
timestamp 28801
transform 1 0 9844 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 28801
transform 1 0 828 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_11
timestamp 28801
transform 1 0 1564 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_39
timestamp 28801
transform 1 0 4140 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_60
timestamp 28801
transform 1 0 6072 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_68
timestamp 28801
transform 1 0 6808 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_97
timestamp 28801
transform 1 0 9476 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_101
timestamp 28801
transform 1 0 9844 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 28801
transform 1 0 828 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_52
timestamp 28801
transform 1 0 5336 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_81
timestamp 28801
transform 1 0 8004 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_85
timestamp 28801
transform 1 0 8372 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_96
timestamp 28801
transform 1 0 9384 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 28801
transform 1 0 828 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_20
timestamp 28801
transform 1 0 2392 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_26
timestamp 28801
transform 1 0 2944 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_34
timestamp 28801
transform 1 0 3680 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_73
timestamp 28801
transform 1 0 7268 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_81
timestamp 28801
transform 1 0 8004 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_96
timestamp 28801
transform 1 0 9384 0 -1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636997256
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_15
timestamp 28801
transform 1 0 1932 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 28801
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_32
timestamp 1636997256
transform 1 0 3496 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_44
timestamp 28801
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_71
timestamp 1636997256
transform 1 0 7084 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 28801
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_93
timestamp 28801
transform 1 0 9108 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_101
timestamp 28801
transform 1 0 9844 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 28801
transform 1 0 828 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_11
timestamp 28801
transform 1 0 1564 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_30
timestamp 28801
transform 1 0 3312 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_38
timestamp 28801
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 28801
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 28801
transform 1 0 828 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_36
timestamp 28801
transform 1 0 3864 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_40
timestamp 28801
transform 1 0 4232 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_61
timestamp 28801
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_79
timestamp 28801
transform 1 0 7820 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 28801
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_101
timestamp 28801
transform 1 0 9844 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_27
timestamp 28801
transform 1 0 3036 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_49
timestamp 28801
transform 1 0 5060 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 28801
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1636997256
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_69
timestamp 28801
transform 1 0 6900 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_73
timestamp 28801
transform 1 0 7268 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_19
timestamp 28801
transform 1 0 2300 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 28801
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_53
timestamp 28801
transform 1 0 5428 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_62
timestamp 28801
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 28801
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 28801
transform 1 0 8372 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636997256
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_15
timestamp 28801
transform 1 0 1932 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_38
timestamp 1636997256
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_50
timestamp 28801
transform 1 0 5152 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_73
timestamp 28801
transform 1 0 7268 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_6
timestamp 28801
transform 1 0 1104 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 28801
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_45
timestamp 28801
transform 1 0 4692 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_62
timestamp 28801
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_101
timestamp 28801
transform 1 0 9844 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_30
timestamp 28801
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_101
timestamp 28801
transform 1 0 9844 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_19
timestamp 28801
transform 1 0 2300 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_51
timestamp 28801
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_74
timestamp 28801
transform 1 0 7360 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 28801
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_101
timestamp 28801
transform 1 0 9844 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 28801
transform -1 0 9476 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 28801
transform 1 0 2392 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 28801
transform 1 0 3496 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 28801
transform 1 0 828 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 28801
transform 1 0 920 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 28801
transform 1 0 7452 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 28801
transform -1 0 9936 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 28801
transform -1 0 9936 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 28801
transform -1 0 5428 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 28801
transform 1 0 6348 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 28801
transform -1 0 3036 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 28801
transform -1 0 9568 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 28801
transform 1 0 4876 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 28801
transform -1 0 9108 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 28801
transform -1 0 9476 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 28801
transform -1 0 7176 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 28801
transform -1 0 1564 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 28801
transform 1 0 3036 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 28801
transform -1 0 3496 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 28801
transform 1 0 3496 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 28801
transform 1 0 5796 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 28801
transform 1 0 5428 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 28801
transform 1 0 7084 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 28801
transform -1 0 6348 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 28801
transform -1 0 8188 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 28801
transform -1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 28801
transform -1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 28801
transform -1 0 9936 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 28801
transform 1 0 9476 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_17
timestamp 28801
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 28801
transform -1 0 10212 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_18
timestamp 28801
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 28801
transform -1 0 10212 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_19
timestamp 28801
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 28801
transform -1 0 10212 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_20
timestamp 28801
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 28801
transform -1 0 10212 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_21
timestamp 28801
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 28801
transform -1 0 10212 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_22
timestamp 28801
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 28801
transform -1 0 10212 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_23
timestamp 28801
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 28801
transform -1 0 10212 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_24
timestamp 28801
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 28801
transform -1 0 10212 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_25
timestamp 28801
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 28801
transform -1 0 10212 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_26
timestamp 28801
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 28801
transform -1 0 10212 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_27
timestamp 28801
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 28801
transform -1 0 10212 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_28
timestamp 28801
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 28801
transform -1 0 10212 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_29
timestamp 28801
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 28801
transform -1 0 10212 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_30
timestamp 28801
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 28801
transform -1 0 10212 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_31
timestamp 28801
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 28801
transform -1 0 10212 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_32
timestamp 28801
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 28801
transform -1 0 10212 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_33
timestamp 28801
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 28801
transform -1 0 10212 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp 28801
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp 28801
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp 28801
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_37
timestamp 28801
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_38
timestamp 28801
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_39
timestamp 28801
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_40
timestamp 28801
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_41
timestamp 28801
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_42
timestamp 28801
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_43
timestamp 28801
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_44
timestamp 28801
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_45
timestamp 28801
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_46
timestamp 28801
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_47
timestamp 28801
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_48
timestamp 28801
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_49
timestamp 28801
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_50
timestamp 28801
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_51
timestamp 28801
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_52
timestamp 28801
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_53
timestamp 28801
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_54
timestamp 28801
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_55
timestamp 28801
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_56
timestamp 28801
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_57
timestamp 28801
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_58
timestamp 28801
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_59
timestamp 28801
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_60
timestamp 28801
transform 1 0 5704 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_61
timestamp 28801
transform 1 0 8280 0 1 9248
box -38 -48 130 592
<< labels >>
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 CLK
port 0 nsew signal input
flabel metal2 s 9494 9957 9550 10757 0 FreeSans 224 90 0 0 CLK_OUT
port 1 nsew signal output
flabel metal2 s 10322 9957 10378 10757 0 FreeSans 224 90 0 0 CLK_OUTn
port 2 nsew signal output
flabel metal2 s 1214 9957 1270 10757 0 FreeSans 224 90 0 0 N[0]
port 3 nsew signal input
flabel metal2 s 2042 9957 2098 10757 0 FreeSans 224 90 0 0 N[1]
port 4 nsew signal input
flabel metal2 s 2870 9957 2926 10757 0 FreeSans 224 90 0 0 N[2]
port 5 nsew signal input
flabel metal2 s 3698 9957 3754 10757 0 FreeSans 224 90 0 0 N[3]
port 6 nsew signal input
flabel metal2 s 4526 9957 4582 10757 0 FreeSans 224 90 0 0 N[4]
port 7 nsew signal input
flabel metal2 s 5354 9957 5410 10757 0 FreeSans 224 90 0 0 N[5]
port 8 nsew signal input
flabel metal2 s 6182 9957 6238 10757 0 FreeSans 224 90 0 0 N[6]
port 9 nsew signal input
flabel metal2 s 7010 9957 7066 10757 0 FreeSans 224 90 0 0 N[7]
port 10 nsew signal input
flabel metal2 s 7838 9957 7894 10757 0 FreeSans 224 90 0 0 N[8]
port 11 nsew signal input
flabel metal2 s 8666 9957 8722 10757 0 FreeSans 224 90 0 0 N[9]
port 12 nsew signal input
flabel metal2 s 386 9957 442 10757 0 FreeSans 224 90 0 0 RESETn
port 13 nsew signal input
flabel metal4 s 4316 496 4636 9840 0 FreeSans 1920 90 0 0 VGND
port 14 nsew ground bidirectional
flabel metal4 s 3656 496 3976 9840 0 FreeSans 1920 90 0 0 VPWR
port 15 nsew power bidirectional
rlabel metal1 5382 9248 5382 9248 0 VGND
rlabel metal1 5382 9792 5382 9792 0 VPWR
rlabel metal1 5106 5066 5106 5066 0 CLK
rlabel metal1 9660 6698 9660 6698 0 CLK_OUT
rlabel metal1 10028 9146 10028 9146 0 CLK_OUTn
rlabel metal1 1288 8398 1288 8398 0 N[0]
rlabel metal1 2070 9044 2070 9044 0 N[1]
rlabel metal1 3082 9486 3082 9486 0 N[2]
rlabel metal1 3634 9486 3634 9486 0 N[3]
rlabel metal1 6026 9588 6026 9588 0 N[4]
rlabel metal1 5520 9486 5520 9486 0 N[5]
rlabel metal1 7314 9554 7314 9554 0 N[6]
rlabel metal1 6118 9520 6118 9520 0 N[7]
rlabel metal1 7958 7276 7958 7276 0 N[8]
rlabel metal2 6578 9044 6578 9044 0 N[9]
rlabel metal1 644 8398 644 8398 0 RESETn
rlabel metal1 7948 5746 7948 5746 0 _000_
rlabel metal1 8224 6222 8224 6222 0 _001_
rlabel metal1 5581 6154 5581 6154 0 _002_
rlabel metal1 2714 3944 2714 3944 0 _003_
rlabel metal2 2162 3706 2162 3706 0 _004_
rlabel via1 3537 2890 3537 2890 0 _005_
rlabel metal1 5101 3638 5101 3638 0 _006_
rlabel metal1 4416 1530 4416 1530 0 _007_
rlabel metal2 6762 1598 6762 1598 0 _008_
rlabel via1 7585 1394 7585 1394 0 _009_
rlabel metal1 8321 2550 8321 2550 0 _010_
rlabel metal1 8592 2958 8592 2958 0 _011_
rlabel via2 4002 3621 4002 3621 0 _012_
rlabel metal1 6210 4080 6210 4080 0 _013_
rlabel metal2 6210 4148 6210 4148 0 _014_
rlabel metal2 6026 5916 6026 5916 0 _015_
rlabel metal1 7820 1870 7820 1870 0 _016_
rlabel metal1 7360 4250 7360 4250 0 _017_
rlabel metal1 6900 4522 6900 4522 0 _018_
rlabel metal1 7130 6222 7130 6222 0 _019_
rlabel metal1 7406 6154 7406 6154 0 _020_
rlabel metal1 7222 4794 7222 4794 0 _021_
rlabel metal1 7176 6154 7176 6154 0 _022_
rlabel metal2 6946 5576 6946 5576 0 _023_
rlabel metal1 6348 4046 6348 4046 0 _024_
rlabel metal1 5704 4046 5704 4046 0 _025_
rlabel metal1 6118 4454 6118 4454 0 _026_
rlabel metal2 4186 5270 4186 5270 0 _027_
rlabel metal1 3818 4114 3818 4114 0 _028_
rlabel metal1 3956 4590 3956 4590 0 _029_
rlabel metal1 4876 4794 4876 4794 0 _030_
rlabel metal1 5566 4794 5566 4794 0 _031_
rlabel metal1 5566 1462 5566 1462 0 _032_
rlabel metal1 6900 5814 6900 5814 0 _033_
rlabel metal1 7218 5882 7218 5882 0 _034_
rlabel metal2 2898 4352 2898 4352 0 _035_
rlabel metal1 2438 3672 2438 3672 0 _036_
rlabel metal2 2346 4182 2346 4182 0 _037_
rlabel metal1 2195 3706 2195 3706 0 _038_
rlabel metal1 5290 2482 5290 2482 0 _039_
rlabel metal1 3726 2312 3726 2312 0 _040_
rlabel metal1 3434 2550 3434 2550 0 _041_
rlabel metal2 7498 4318 7498 4318 0 _042_
rlabel metal1 5796 1870 5796 1870 0 _043_
rlabel metal1 5152 1190 5152 1190 0 _044_
rlabel via1 4730 1530 4730 1530 0 _045_
rlabel metal1 6440 2074 6440 2074 0 _046_
rlabel metal2 8050 2142 8050 2142 0 _047_
rlabel metal1 6762 1870 6762 1870 0 _048_
rlabel metal1 7130 1836 7130 1836 0 _049_
rlabel metal1 7314 2312 7314 2312 0 _050_
rlabel metal1 7866 2856 7866 2856 0 _051_
rlabel metal1 8188 2074 8188 2074 0 _052_
rlabel metal1 7406 3162 7406 3162 0 _053_
rlabel metal1 7406 7820 7406 7820 0 clknet_0_CLK
rlabel metal1 966 4692 966 4692 0 clknet_2_0__leaf_CLK
rlabel metal1 8188 2482 8188 2482 0 clknet_2_1__leaf_CLK
rlabel metal2 2254 6494 2254 6494 0 clknet_2_2__leaf_CLK
rlabel metal1 7314 9044 7314 9044 0 clknet_2_3__leaf_CLK
rlabel metal1 3542 6324 3542 6324 0 counter\[0\]
rlabel metal1 2530 4624 2530 4624 0 counter\[1\]
rlabel metal2 2622 3740 2622 3740 0 counter\[2\]
rlabel metal1 2714 3468 2714 3468 0 counter\[3\]
rlabel via2 6118 4029 6118 4029 0 counter\[4\]
rlabel metal1 5106 2448 5106 2448 0 counter\[5\]
rlabel metal1 6302 2618 6302 2618 0 counter\[6\]
rlabel metal1 7912 1802 7912 1802 0 counter\[7\]
rlabel metal2 8050 3638 8050 3638 0 counter\[8\]
rlabel metal1 9614 1938 9614 1938 0 counter\[9\]
rlabel metal1 690 9010 690 9010 0 n0\[0\]
rlabel metal1 690 6630 690 6630 0 n0\[1\]
rlabel metal1 5290 7412 5290 7412 0 n0\[2\]
rlabel metal2 1610 9316 1610 9316 0 n0\[3\]
rlabel metal2 3634 9146 3634 9146 0 n0\[4\]
rlabel metal1 6026 9146 6026 9146 0 n0\[5\]
rlabel metal1 7360 9146 7360 9146 0 n0\[6\]
rlabel metal1 9246 7922 9246 7922 0 n0\[7\]
rlabel metal2 9798 8772 9798 8772 0 n0\[8\]
rlabel metal1 9752 5746 9752 5746 0 n0\[9\]
rlabel metal1 3220 6222 3220 6222 0 n\[0\]
rlabel metal2 3266 5372 3266 5372 0 n\[1\]
rlabel metal1 4830 4726 4830 4726 0 n\[2\]
rlabel metal1 4048 4726 4048 4726 0 n\[3\]
rlabel metal1 6348 4658 6348 4658 0 n\[4\]
rlabel metal2 6026 7514 6026 7514 0 n\[5\]
rlabel metal2 6578 6698 6578 6698 0 n\[6\]
rlabel metal2 7774 5644 7774 5644 0 n\[7\]
rlabel metal1 8648 4046 8648 4046 0 n\[8\]
rlabel metal1 8832 4658 8832 4658 0 n\[9\]
rlabel metal1 1656 8602 1656 8602 0 net1
rlabel metal1 7176 8602 7176 8602 0 net10
rlabel via1 1145 7310 1145 7310 0 net11
rlabel metal2 9890 6630 9890 6630 0 net12
rlabel metal2 9154 7446 9154 7446 0 net13
rlabel via1 7125 8330 7125 8330 0 net14
rlabel metal1 3296 8330 3296 8330 0 net15
rlabel metal1 5004 8398 5004 8398 0 net16
rlabel metal1 1686 8330 1686 8330 0 net17
rlabel metal1 1778 6154 1778 6154 0 net18
rlabel metal1 7692 7310 7692 7310 0 net19
rlabel metal2 2806 7820 2806 7820 0 net2
rlabel metal1 9384 5882 9384 5882 0 net20
rlabel metal1 8893 6902 8893 6902 0 net21
rlabel metal1 4319 6834 4319 6834 0 net22
rlabel metal1 7002 7922 7002 7922 0 net23
rlabel metal1 2249 5814 2249 5814 0 net24
rlabel metal1 8234 6086 8234 6086 0 net25
rlabel metal1 5704 5882 5704 5882 0 net26
rlabel metal2 7038 5610 7038 5610 0 net27
rlabel metal1 7590 2992 7590 2992 0 net28
rlabel metal1 6256 3570 6256 3570 0 net29
rlabel metal1 3440 7310 3440 7310 0 net3
rlabel metal2 3542 9214 3542 9214 0 net4
rlabel metal1 5397 9418 5397 9418 0 net5
rlabel metal1 5009 9078 5009 9078 0 net6
rlabel metal1 6619 9010 6619 9010 0 net7
rlabel metal1 7493 9078 7493 9078 0 net8
rlabel metal2 8142 7922 8142 7922 0 net9
rlabel metal1 5842 5610 5842 5610 0 resetn
rlabel metal2 2898 7004 2898 7004 0 resetn0
<< properties >>
string FIXED_BBOX 0 0 10773 10757
<< end >>
