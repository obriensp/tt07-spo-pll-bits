* testing extracted vco

V1 vdd GND {VDD}
V2 vss GND 0

* frequency control voltage (higher voltage = higher frequency)
V3 vcont GND {VCONT}

* digital signals for vco's capacitive loads (high = more load, slower frequency)
V4 s0 GND {S0}
V5 s1 GND {S1}

*.subckt vco_parax s0 s1 out vcont vss vdd
x1 s0 s1 out vcont vss net_measured_vdd vco_parax

* measure current consumed by vco
Vmeas vdd net_measured_vdd 0
.save i(vmeas)

.include vco_prefix.spice
.include ../mag/vco.sim.spice

*.option savecurrents
.control
  save all
  tran 10p 500n 100n
  wrdata out/vco_current.txt vmeas#branch
  linearize
  fft v(out)
  wrdata out/vco_fft.txt mag(V(out))
  quit
.endc

.global GND
.end
