magic
tech sky130A
magscale 1 2
timestamp 1717212334
<< pwell >>
rect 1330 -2580 1490 -2090
<< viali >>
rect 1852 -1362 2010 -1328
rect 2272 -1362 2430 -1328
rect 1432 -2604 1590 -2570
rect 1852 -2604 2010 -2570
rect 2272 -2604 2430 -2570
<< metal1 >>
rect 1040 -1328 2570 -1220
rect 1040 -1362 1852 -1328
rect 2010 -1362 2272 -1328
rect 2430 -1362 2570 -1328
rect 1040 -1370 2570 -1362
rect 1040 -1420 1240 -1370
rect 1040 -1594 1240 -1520
rect 1278 -1594 1284 -1593
rect 1040 -1645 1284 -1594
rect 1336 -1645 1342 -1593
rect 1780 -1630 1910 -1370
rect 1950 -1494 2090 -1450
rect 1950 -1546 2025 -1494
rect 2077 -1546 2090 -1494
rect 1950 -1630 2090 -1546
rect 2200 -1630 2330 -1370
rect 2370 -1630 2510 -1450
rect 2640 -1591 2840 -1520
rect 1040 -1720 1240 -1645
rect 2050 -1680 2090 -1630
rect 1870 -1760 1880 -1680
rect 1960 -1760 1970 -1680
rect 2050 -1740 2380 -1680
rect 1040 -1914 1240 -1830
rect 1040 -1946 1526 -1914
rect 1040 -2030 1240 -1946
rect 1494 -2000 1526 -1946
rect 1470 -2060 1550 -2000
rect 1870 -2060 1880 -1970
rect 1970 -2060 1980 -1970
rect 1040 -2230 1240 -2170
rect 1040 -2310 1270 -2230
rect 1340 -2310 1350 -2230
rect 1040 -2370 1240 -2310
rect 1040 -2500 1240 -2450
rect 1380 -2500 1490 -2090
rect 1530 -2110 1910 -2090
rect 2050 -2100 2090 -1740
rect 2470 -1780 2510 -1630
rect 2555 -1649 2561 -1591
rect 2619 -1649 2840 -1591
rect 2640 -1720 2840 -1649
rect 2440 -1860 2450 -1780
rect 2530 -1860 2540 -1780
rect 2300 -2060 2310 -1970
rect 2400 -2060 2410 -1970
rect 1530 -2470 1760 -2110
rect 1850 -2470 1910 -2110
rect 1950 -2460 2090 -2100
rect 2160 -2110 2330 -2090
rect 2470 -2100 2510 -1860
rect 1530 -2490 1910 -2470
rect 2160 -2470 2180 -2110
rect 2270 -2470 2330 -2110
rect 2370 -2241 2510 -2100
rect 2640 -2241 2840 -2170
rect 2370 -2299 2840 -2241
rect 2370 -2460 2510 -2299
rect 2640 -2370 2840 -2299
rect 2160 -2490 2330 -2470
rect 1040 -2560 1490 -2500
rect 1040 -2570 2570 -2560
rect 1040 -2604 1432 -2570
rect 1590 -2604 1852 -2570
rect 2010 -2604 2272 -2570
rect 2430 -2604 2570 -2570
rect 1040 -2650 2570 -2604
<< via1 >>
rect 1284 -1645 1336 -1593
rect 2025 -1546 2077 -1494
rect 1880 -1760 1960 -1680
rect 1880 -2060 1970 -1970
rect 1270 -2310 1340 -2230
rect 2561 -1649 2619 -1591
rect 2450 -1860 2530 -1780
rect 2310 -2060 2400 -1970
rect 1760 -2470 1850 -2110
rect 2180 -2470 2270 -2110
<< metal2 >>
rect 2025 -1494 2077 -1488
rect 2025 -1552 2077 -1546
rect 1284 -1593 1336 -1587
rect 2029 -1598 2072 -1552
rect 2561 -1591 2619 -1585
rect 1336 -1635 1646 -1602
rect 1284 -1651 1336 -1645
rect 1613 -1893 1646 -1635
rect 2029 -1641 2561 -1598
rect 2561 -1655 2619 -1649
rect 1880 -1680 1960 -1670
rect 1880 -1770 1960 -1760
rect 1890 -1800 1940 -1770
rect 2450 -1780 2530 -1770
rect 1890 -1850 2450 -1800
rect 2450 -1870 2530 -1860
rect 1613 -1926 2366 -1893
rect 2333 -1960 2366 -1926
rect 1880 -1970 1970 -1960
rect 1296 -2025 1880 -1996
rect 1296 -2220 1325 -2025
rect 1880 -2070 1970 -2060
rect 2310 -1970 2400 -1960
rect 2310 -2070 2400 -2060
rect 1760 -2110 1850 -2100
rect 2180 -2110 2270 -2100
rect 1270 -2230 1340 -2220
rect 1270 -2320 1340 -2310
rect 1850 -2470 2180 -2110
rect 1760 -2480 1850 -2470
rect 2180 -2480 2270 -2470
use sky130_fd_pr__nfet_01v8_26NUYT  sky130_fd_pr__nfet_01v8_26NUYT_0
timestamp 1717210983
transform 1 0 2351 0 1 -2261
box -211 -379 211 379
use sky130_fd_pr__pfet_01v8_7PK3FC  sky130_fd_pr__pfet_01v8_7PK3FC_0
timestamp 1717210983
transform 1 0 2351 0 1 -1576
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_26NUYT  XM1
timestamp 1717210983
transform 1 0 1931 0 1 -2261
box -211 -379 211 379
use sky130_fd_pr__nfet_01v8_26NUYT  XM4
timestamp 1717210983
transform 1 0 1511 0 1 -2261
box -211 -379 211 379
use sky130_fd_pr__pfet_01v8_7PK3FC  XM11
timestamp 1717210983
transform 1 0 1931 0 1 -1576
box -211 -284 211 284
<< labels >>
flabel metal1 1040 -2370 1240 -2170 0 FreeSans 256 0 0 0 d_n
port 5 nsew
flabel metal1 1040 -1720 1240 -1520 0 FreeSans 256 0 0 0 d
port 4 nsew
flabel metal1 1040 -2030 1240 -1830 0 FreeSans 256 0 0 0 clk
port 6 nsew
flabel metal1 1040 -2650 1240 -2450 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 1040 -1420 1240 -1220 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 2640 -1720 2840 -1520 0 FreeSans 256 0 0 0 q
port 3 nsew
flabel metal1 2640 -2370 2840 -2170 0 FreeSans 256 0 0 0 q_n
port 2 nsew
<< end >>
