magic
tech sky130A
magscale 1 2
timestamp 1716529149
<< metal1 >>
rect 16182 15182 16192 15382
rect 16392 15182 16402 15382
rect 16508 15182 16518 15382
rect 16718 15182 16728 15382
rect 16822 15182 16832 15382
rect 17032 15182 17042 15382
rect 15528 14066 15538 14270
rect 15762 14066 15772 14270
rect 15154 13558 15164 13758
rect 15364 13558 15374 13758
rect 15826 13560 15836 13760
rect 16036 13560 16046 13760
rect 16184 13344 16194 13544
rect 16394 13344 16404 13544
rect 16520 13444 16720 13650
rect 17144 13558 17154 13758
rect 17354 13558 17364 13758
rect 17542 13558 17552 13758
rect 17752 13558 17762 13758
rect 16824 13344 16834 13544
rect 17034 13344 17044 13544
rect 15530 12228 15540 12432
rect 15764 12228 15774 12432
rect 15156 11720 15166 11920
rect 15366 11720 15376 11920
rect 15828 11722 15838 11922
rect 16038 11722 16048 11922
rect 16188 11500 16198 11700
rect 16398 11500 16408 11700
rect 16522 11670 16722 11876
rect 17146 11720 17156 11920
rect 17356 11720 17366 11920
rect 17544 11720 17554 11920
rect 17754 11720 17764 11920
rect 16828 11500 16838 11700
rect 17038 11500 17048 11700
rect 15534 10384 15544 10588
rect 15768 10384 15778 10588
rect 15160 9876 15170 10076
rect 15370 9876 15380 10076
rect 15832 9878 15842 10078
rect 16042 9878 16052 10078
rect 16516 9874 16526 10074
rect 16726 9874 16736 10074
rect 17150 9876 17160 10076
rect 17360 9876 17370 10076
rect 17548 9876 17558 10076
rect 17758 9876 17768 10076
<< via1 >>
rect 16192 15182 16392 15382
rect 16518 15182 16718 15382
rect 16832 15182 17032 15382
rect 15538 14066 15762 14270
rect 15164 13558 15364 13758
rect 15836 13560 16036 13760
rect 16194 13344 16394 13544
rect 17154 13558 17354 13758
rect 17552 13558 17752 13758
rect 16834 13344 17034 13544
rect 15540 12228 15764 12432
rect 15166 11720 15366 11920
rect 15838 11722 16038 11922
rect 16198 11500 16398 11700
rect 17156 11720 17356 11920
rect 17554 11720 17754 11920
rect 16838 11500 17038 11700
rect 15544 10384 15768 10588
rect 15170 9876 15370 10076
rect 15842 9878 16042 10078
rect 16526 9874 16726 10074
rect 17160 9876 17360 10076
rect 17558 9876 17758 10076
<< metal2 >>
rect 16192 15382 16392 15392
rect 16192 15172 16392 15182
rect 16518 15382 16718 15392
rect 16518 15172 16718 15182
rect 16832 15382 17032 15392
rect 16832 15172 17032 15182
rect 15538 14270 15762 14280
rect 15204 13768 15332 14134
rect 15538 14056 15762 14066
rect 15164 13758 15364 13768
rect 15164 13548 15364 13558
rect 15204 11930 15332 13548
rect 15584 12442 15712 14056
rect 15836 13760 16036 13770
rect 15836 13550 16036 13560
rect 16238 13554 16366 15172
rect 16864 13554 16992 15172
rect 17590 13768 17718 14146
rect 17154 13758 17354 13768
rect 15540 12432 15764 12442
rect 15540 12218 15764 12228
rect 15166 11920 15366 11930
rect 15166 11710 15366 11720
rect 15204 10086 15332 11710
rect 15584 10598 15712 12218
rect 15876 11932 16004 13550
rect 16194 13544 16394 13554
rect 16194 13334 16394 13344
rect 16834 13544 17034 13554
rect 17154 13548 17354 13558
rect 17552 13758 17752 13768
rect 17552 13548 17752 13558
rect 16834 13334 17034 13344
rect 15838 11922 16038 11932
rect 15838 11712 16038 11722
rect 15544 10588 15768 10598
rect 15544 10374 15584 10384
rect 15712 10374 15768 10384
rect 15876 10088 16004 11712
rect 16238 11710 16366 13334
rect 16864 11710 16992 13334
rect 17194 11930 17322 13548
rect 17590 11930 17718 13548
rect 17156 11920 17356 11930
rect 17156 11710 17356 11720
rect 17554 11920 17754 11930
rect 17554 11710 17754 11720
rect 16198 11700 16398 11710
rect 16198 11490 16238 11500
rect 16366 11490 16398 11500
rect 16838 11700 17038 11710
rect 16838 11490 17038 11500
rect 15170 10076 15370 10086
rect 15170 9866 15204 9876
rect 15332 9866 15370 9876
rect 15842 10078 16042 10088
rect 17194 10086 17322 11710
rect 17590 10086 17718 11710
rect 15842 9868 15876 9878
rect 16004 9868 16042 9878
rect 16526 10074 16726 10084
rect 16526 9864 16567 9874
rect 16669 9864 16726 9874
rect 17160 10076 17360 10086
rect 17160 9866 17194 9876
rect 17322 9866 17360 9876
rect 17558 10076 17758 10086
rect 17558 9866 17590 9876
rect 17718 9866 17758 9876
<< via2 >>
rect 16518 15182 16718 15382
rect 16526 9874 16726 10074
<< metal3 >>
rect 16508 15382 16728 15387
rect 16508 15182 16518 15382
rect 16718 15182 16728 15382
rect 16508 15177 16728 15182
rect 16567 10079 16669 15177
rect 16516 10074 16736 10079
rect 16516 9874 16526 10074
rect 16726 9874 16736 10074
rect 16516 9869 16736 9874
rect 16528 9868 16734 9869
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 1000 500 44152
rect 9800 1000 10100 44152
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 200
use delay_stage  delay_stage_0 ~/Development/spo/vlsi/tt07-spo-pll/mag
timestamp 1716529149
transform 1 0 14706 0 1 15462
box 208 -1906 3270 -80
use delay_stage  delay_stage_1
timestamp 1716529149
transform 1 0 14712 0 1 11780
box 208 -1906 3270 -80
use delay_stage  delay_stage_2
timestamp 1716529149
transform 1 0 14708 0 1 13624
box 208 -1906 3270 -80
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
