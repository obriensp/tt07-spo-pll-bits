magic
tech sky130A
magscale 1 2
timestamp 1717172438
<< metal3 >>
rect 29494 26732 29570 26738
rect 28472 26668 28478 26732
rect 28542 26730 28548 26732
rect 29494 26730 29500 26732
rect 28542 26670 29500 26730
rect 28542 26668 28548 26670
rect 29494 26668 29500 26670
rect 29564 26668 29570 26732
rect 29494 26662 29570 26668
rect 190 9249 510 9260
rect 190 8951 201 9249
rect 499 9212 510 9249
rect 499 8989 15061 9212
rect 499 8951 510 8989
rect 190 8940 510 8951
rect 9801 8679 10099 8685
rect 10099 8429 14591 8631
rect 14838 8429 15061 8989
rect 15302 9187 31446 9188
rect 15302 9052 31310 9187
rect 31445 9052 31451 9187
rect 15302 9051 31446 9052
rect 15302 8412 15439 9051
rect 15680 8480 15690 8610
rect 15820 8480 15830 8610
rect 16080 8480 16090 8610
rect 16220 8480 16230 8610
rect 16480 8480 16490 8610
rect 16620 8480 16630 8610
rect 9801 8375 10099 8381
<< via3 >>
rect 28478 26668 28542 26732
rect 29500 26668 29564 26732
rect 201 8951 499 9249
rect 9801 8381 10099 8679
rect 31310 9052 31445 9187
rect 15690 8480 15820 8610
rect 16090 8480 16220 8610
rect 16490 8480 16620 8610
<< metal4 >>
rect 798 44460 858 45152
rect 1534 44800 1594 45152
rect 2270 44800 2330 45152
rect 3006 44800 3066 45152
rect 3742 44800 3802 45152
rect 4478 44800 4538 45152
rect 5214 44800 5274 45152
rect 5950 44800 6010 45152
rect 6686 44800 6746 45152
rect 7422 44800 7482 45152
rect 8158 44800 8218 45152
rect 8894 44800 8954 45152
rect 9630 44800 9690 45152
rect 10366 44800 10426 45152
rect 11102 44800 11162 45152
rect 11838 44800 11898 45152
rect 12574 44800 12634 45152
rect 13310 44800 13370 45152
rect 14046 44800 14106 45152
rect 14782 44800 14842 45152
rect 15518 44800 15578 45152
rect 16254 44800 16314 45152
rect 16990 44800 17050 45152
rect 1220 44460 17270 44800
rect 798 44400 17270 44460
rect 200 9249 500 44152
rect 1220 44110 17270 44400
rect 200 8951 201 9249
rect 499 8951 500 9249
rect 200 5431 500 8951
rect 9800 8679 10100 44110
rect 17726 13650 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28477 26732 28543 26733
rect 28477 26668 28478 26732
rect 28542 26668 28543 26732
rect 28477 26667 28543 26668
rect 15720 13590 17786 13650
rect 15720 8840 15780 13590
rect 28480 10400 28540 26667
rect 16110 10340 28540 10400
rect 16110 8840 16170 10340
rect 28766 10040 28826 45152
rect 29502 26733 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 29499 26732 29565 26733
rect 29499 26668 29500 26732
rect 29564 26668 29565 26732
rect 29499 26667 29565 26668
rect 16510 9980 28826 10040
rect 16510 8840 16570 9980
rect 28766 9960 28826 9980
rect 31309 9187 31446 9188
rect 31309 9052 31310 9187
rect 31445 9052 31446 9187
rect 9800 8381 9801 8679
rect 10099 8381 10100 8679
rect 15690 8611 15820 8840
rect 16090 8611 16220 8840
rect 16490 8611 16620 8840
rect 15689 8610 15821 8611
rect 15689 8480 15690 8610
rect 15820 8480 15821 8610
rect 15689 8479 15821 8480
rect 16089 8610 16221 8611
rect 16089 8480 16090 8610
rect 16220 8480 16221 8610
rect 16089 8479 16221 8480
rect 16489 8610 16621 8611
rect 16489 8480 16490 8610
rect 16620 8480 16621 8610
rect 16489 8479 16621 8480
rect 15690 8475 15820 8479
rect 199 5139 501 5431
rect 200 1000 500 5139
rect 9800 2951 10100 8381
rect 9799 2659 10101 2951
rect 9800 1000 10100 2659
rect 31309 200 31446 9052
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 200
use vco  vco_0
timestamp 1717119155
transform 1 0 15000 0 1 6406
box -530 -1206 4600 2230
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 0 FreeSans 1600 0 0 0 VPWR
port 52 nsew
flabel space 9801 1000 10101 44152 0 FreeSans 1600 0 0 0 VGND
port 51 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
