MACRO tt_um_obriensp_pll
  CLASS BLOCK ;
  FOREIGN tt_um_obriensp_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.650000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.350000 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 27.913649 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 25.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 13.300 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 94.885 42.535 95.055 42.725 ;
        RECT 85.545 42.285 90.640 42.535 ;
        RECT 93.435 42.365 95.195 42.535 ;
        RECT 92.940 42.320 95.195 42.365 ;
        RECT 92.000 42.285 95.195 42.320 ;
        RECT 85.545 41.855 95.195 42.285 ;
        RECT 85.545 41.625 87.565 41.855 ;
        RECT 86.645 41.605 87.565 41.625 ;
        RECT 90.640 41.685 93.870 41.855 ;
        RECT 90.640 41.640 92.930 41.685 ;
        RECT 95.215 41.665 95.645 42.450 ;
        RECT 90.640 41.605 91.990 41.640 ;
      LAYER nwell ;
        RECT 85.350 39.730 95.850 41.335 ;
        RECT 75.000 37.170 97.950 38.330 ;
        RECT 72.750 33.330 97.950 37.170 ;
        RECT 75.000 31.130 97.950 33.330 ;
      LAYER pwell ;
        RECT 75.000 30.720 97.950 31.080 ;
        RECT 72.750 26.930 97.950 30.720 ;
        RECT 75.000 26.030 97.950 26.930 ;
      LAYER li1 ;
        RECT 85.540 42.555 95.660 42.725 ;
        RECT 85.625 40.175 85.885 42.385 ;
        RECT 86.135 42.095 86.305 42.555 ;
        RECT 86.475 42.215 87.470 42.385 ;
        RECT 88.000 42.225 88.170 42.385 ;
        RECT 86.475 41.925 86.645 42.215 ;
        RECT 87.300 42.055 87.470 42.215 ;
        RECT 87.640 42.055 88.170 42.225 ;
        RECT 86.075 41.755 86.645 41.925 ;
        RECT 86.815 41.875 86.990 42.045 ;
        RECT 86.075 40.975 86.245 41.755 ;
        RECT 86.815 41.715 87.230 41.875 ;
        RECT 86.820 41.705 87.230 41.715 ;
        RECT 86.555 41.365 87.010 41.535 ;
        RECT 86.075 40.805 86.725 40.975 ;
        RECT 87.640 40.885 87.810 42.055 ;
        RECT 88.515 41.985 88.690 42.315 ;
        RECT 88.860 42.175 89.190 42.555 ;
        RECT 87.980 41.705 88.220 41.875 ;
        RECT 86.055 40.005 86.385 40.385 ;
        RECT 86.555 40.345 86.725 40.805 ;
        RECT 87.025 40.655 87.810 40.885 ;
        RECT 87.025 40.515 87.355 40.655 ;
        RECT 88.050 40.505 88.220 41.705 ;
        RECT 88.515 41.535 88.685 41.985 ;
        RECT 89.460 41.925 89.705 42.345 ;
        RECT 89.880 42.095 90.050 42.555 ;
        RECT 90.220 42.215 91.820 42.385 ;
        RECT 90.220 42.175 90.575 42.215 ;
        RECT 90.810 41.925 90.980 42.045 ;
        RECT 89.460 41.755 90.980 41.925 ;
        RECT 90.810 41.715 90.980 41.755 ;
        RECT 91.150 41.795 91.480 42.045 ;
        RECT 91.650 41.845 91.820 42.215 ;
        RECT 92.110 41.835 92.400 42.555 ;
        RECT 93.110 42.215 94.185 42.385 ;
        RECT 91.150 41.720 91.465 41.795 ;
        RECT 88.395 41.365 88.685 41.535 ;
        RECT 87.510 40.345 87.840 40.385 ;
        RECT 86.555 40.175 87.840 40.345 ;
        RECT 88.010 40.175 88.220 40.505 ;
        RECT 88.515 40.505 88.685 41.365 ;
        RECT 88.855 40.965 89.145 41.645 ;
        RECT 89.620 40.965 89.950 41.585 ;
        RECT 90.155 40.965 90.400 41.585 ;
        RECT 90.795 41.535 91.125 41.545 ;
        RECT 90.740 41.375 91.125 41.535 ;
        RECT 90.740 41.365 90.910 41.375 ;
        RECT 91.295 41.195 91.465 41.720 ;
        RECT 90.705 41.025 91.465 41.195 ;
        RECT 89.470 40.555 90.535 40.725 ;
        RECT 88.515 40.175 88.700 40.505 ;
        RECT 88.870 40.005 89.220 40.385 ;
        RECT 89.470 40.175 89.640 40.555 ;
        RECT 89.810 40.005 90.140 40.385 ;
        RECT 90.365 40.345 90.535 40.555 ;
        RECT 90.705 40.515 91.035 41.025 ;
        RECT 91.205 40.345 91.375 40.855 ;
        RECT 91.635 40.645 91.935 41.645 ;
        RECT 92.580 41.535 92.940 42.210 ;
        RECT 93.110 41.880 93.280 42.215 ;
        RECT 93.450 41.875 93.790 42.045 ;
        RECT 93.500 41.705 93.790 41.875 ;
        RECT 94.015 42.005 94.185 42.215 ;
        RECT 94.355 42.175 94.685 42.555 ;
        RECT 94.855 42.005 95.025 42.380 ;
        RECT 94.015 41.835 95.025 42.005 ;
        RECT 95.285 41.830 95.575 42.555 ;
        RECT 92.580 41.355 93.120 41.535 ;
        RECT 92.580 41.245 92.940 41.355 ;
        RECT 92.135 41.015 92.940 41.245 ;
        RECT 93.620 41.185 93.790 41.705 ;
        RECT 93.155 41.015 93.790 41.185 ;
        RECT 93.960 41.025 94.395 41.645 ;
        RECT 94.705 41.025 95.050 41.645 ;
        RECT 90.365 40.175 91.375 40.345 ;
        RECT 91.635 40.005 91.965 40.385 ;
        RECT 92.135 40.175 92.485 41.015 ;
        RECT 92.655 40.345 92.825 40.845 ;
        RECT 93.155 40.685 93.325 41.015 ;
        RECT 92.995 40.515 93.325 40.685 ;
        RECT 93.495 40.675 95.025 40.845 ;
        RECT 93.495 40.515 93.665 40.675 ;
        RECT 94.015 40.345 94.185 40.505 ;
        RECT 92.655 40.175 94.185 40.345 ;
        RECT 94.355 40.005 94.685 40.385 ;
        RECT 94.855 40.175 95.025 40.675 ;
        RECT 95.285 40.005 95.575 41.170 ;
        RECT 85.540 39.835 95.660 40.005 ;
        RECT 74.530 37.800 75.020 38.290 ;
        RECT 75.400 37.920 77.110 38.090 ;
        RECT 77.950 37.920 79.660 38.090 ;
        RECT 80.500 37.920 82.210 38.090 ;
        RECT 83.050 37.920 84.760 38.090 ;
        RECT 85.600 37.920 87.310 38.090 ;
        RECT 88.150 37.920 89.860 38.090 ;
        RECT 90.700 37.920 92.410 38.090 ;
        RECT 93.250 37.920 94.960 38.090 ;
        RECT 95.800 37.920 97.510 38.090 ;
        RECT 72.930 36.820 74.830 36.990 ;
        RECT 72.930 33.680 73.100 36.820 ;
        RECT 73.500 34.410 73.670 36.450 ;
        RECT 74.090 34.410 74.260 36.450 ;
        RECT 73.715 34.025 74.045 34.195 ;
        RECT 74.660 33.680 74.830 36.820 ;
        RECT 75.800 35.510 75.970 37.550 ;
        RECT 76.540 35.510 76.710 37.550 ;
        RECT 76.030 35.125 76.480 35.295 ;
        RECT 77.110 35.015 77.280 37.685 ;
        RECT 78.350 35.510 78.520 37.550 ;
        RECT 79.090 35.510 79.260 37.550 ;
        RECT 78.580 35.125 79.030 35.295 ;
        RECT 79.660 35.015 79.830 37.685 ;
        RECT 80.900 35.510 81.070 37.550 ;
        RECT 81.640 35.510 81.810 37.550 ;
        RECT 81.130 35.125 81.580 35.295 ;
        RECT 82.210 35.015 82.380 37.685 ;
        RECT 83.450 35.510 83.620 37.550 ;
        RECT 84.190 35.510 84.360 37.550 ;
        RECT 83.680 35.125 84.130 35.295 ;
        RECT 84.760 35.015 84.930 37.685 ;
        RECT 86.000 35.510 86.170 37.550 ;
        RECT 86.740 35.510 86.910 37.550 ;
        RECT 86.230 35.125 86.680 35.295 ;
        RECT 87.310 35.015 87.480 37.685 ;
        RECT 88.550 35.510 88.720 37.550 ;
        RECT 89.290 35.510 89.460 37.550 ;
        RECT 88.780 35.125 89.230 35.295 ;
        RECT 89.860 35.015 90.030 37.685 ;
        RECT 91.100 35.510 91.270 37.550 ;
        RECT 91.840 35.510 92.010 37.550 ;
        RECT 91.330 35.125 91.780 35.295 ;
        RECT 92.410 35.015 92.580 37.685 ;
        RECT 93.650 35.510 93.820 37.550 ;
        RECT 94.390 35.510 94.560 37.550 ;
        RECT 93.880 35.125 94.330 35.295 ;
        RECT 94.960 35.015 95.130 37.685 ;
        RECT 96.200 35.510 96.370 37.550 ;
        RECT 96.940 35.510 97.110 37.550 ;
        RECT 96.430 35.125 96.880 35.295 ;
        RECT 97.510 35.015 97.680 37.685 ;
        RECT 72.930 33.510 74.830 33.680 ;
        RECT 75.800 32.210 75.970 34.250 ;
        RECT 76.540 32.210 76.710 34.250 ;
        RECT 78.350 32.210 78.520 34.250 ;
        RECT 79.090 32.210 79.260 34.250 ;
        RECT 80.900 32.210 81.070 34.250 ;
        RECT 81.640 32.210 81.810 34.250 ;
        RECT 83.450 32.210 83.620 34.250 ;
        RECT 84.190 32.210 84.360 34.250 ;
        RECT 86.000 32.210 86.170 34.250 ;
        RECT 86.740 32.210 86.910 34.250 ;
        RECT 88.550 32.210 88.720 34.250 ;
        RECT 89.290 32.210 89.460 34.250 ;
        RECT 91.100 32.210 91.270 34.250 ;
        RECT 91.840 32.210 92.010 34.250 ;
        RECT 93.650 32.210 93.820 34.250 ;
        RECT 94.390 32.210 94.560 34.250 ;
        RECT 96.200 32.210 96.370 34.250 ;
        RECT 96.940 32.210 97.110 34.250 ;
        RECT 76.030 31.825 76.480 31.995 ;
        RECT 78.580 31.825 79.030 31.995 ;
        RECT 81.130 31.825 81.580 31.995 ;
        RECT 83.680 31.825 84.130 31.995 ;
        RECT 86.230 31.825 86.680 31.995 ;
        RECT 88.780 31.825 89.230 31.995 ;
        RECT 91.330 31.825 91.780 31.995 ;
        RECT 93.880 31.825 94.330 31.995 ;
        RECT 96.430 31.825 96.880 31.995 ;
        RECT 75.230 30.720 77.280 30.890 ;
        RECT 72.930 30.370 74.830 30.540 ;
        RECT 72.930 27.280 73.100 30.370 ;
        RECT 73.500 27.960 73.670 30.000 ;
        RECT 74.090 27.960 74.260 30.000 ;
        RECT 73.715 27.620 74.045 27.790 ;
        RECT 74.660 27.280 74.830 30.370 ;
        RECT 72.930 27.110 74.830 27.280 ;
        RECT 75.230 28.640 75.400 30.720 ;
        RECT 76.030 30.210 76.480 30.380 ;
        RECT 75.800 29.000 75.970 30.040 ;
        RECT 76.540 29.000 76.710 30.040 ;
        RECT 77.110 28.640 77.280 30.720 ;
        RECT 75.230 28.460 77.280 28.640 ;
        RECT 72.430 26.060 72.920 26.550 ;
        RECT 75.230 26.380 75.400 28.460 ;
        RECT 76.030 27.960 76.480 28.130 ;
        RECT 75.800 26.750 75.970 27.790 ;
        RECT 76.540 26.750 76.710 27.790 ;
        RECT 77.110 26.380 77.280 28.460 ;
        RECT 75.230 26.210 77.280 26.380 ;
        RECT 77.780 30.720 79.830 30.890 ;
        RECT 77.780 28.640 77.950 30.720 ;
        RECT 78.580 30.210 79.030 30.380 ;
        RECT 78.350 29.000 78.520 30.040 ;
        RECT 79.090 29.000 79.260 30.040 ;
        RECT 79.660 28.640 79.830 30.720 ;
        RECT 77.780 28.460 79.830 28.640 ;
        RECT 77.780 26.380 77.950 28.460 ;
        RECT 78.580 27.960 79.030 28.130 ;
        RECT 78.350 26.750 78.520 27.790 ;
        RECT 79.090 26.750 79.260 27.790 ;
        RECT 79.660 26.380 79.830 28.460 ;
        RECT 77.780 26.210 79.830 26.380 ;
        RECT 80.330 30.720 82.380 30.890 ;
        RECT 80.330 28.640 80.500 30.720 ;
        RECT 81.130 30.210 81.580 30.380 ;
        RECT 80.900 29.000 81.070 30.040 ;
        RECT 81.640 29.000 81.810 30.040 ;
        RECT 82.210 28.640 82.380 30.720 ;
        RECT 80.330 28.460 82.380 28.640 ;
        RECT 80.330 26.380 80.500 28.460 ;
        RECT 81.130 27.960 81.580 28.130 ;
        RECT 80.900 26.750 81.070 27.790 ;
        RECT 81.640 26.750 81.810 27.790 ;
        RECT 82.210 26.380 82.380 28.460 ;
        RECT 80.330 26.210 82.380 26.380 ;
        RECT 82.880 30.720 84.930 30.890 ;
        RECT 82.880 28.640 83.050 30.720 ;
        RECT 83.680 30.210 84.130 30.380 ;
        RECT 83.450 29.000 83.620 30.040 ;
        RECT 84.190 29.000 84.360 30.040 ;
        RECT 84.760 28.640 84.930 30.720 ;
        RECT 82.880 28.460 84.930 28.640 ;
        RECT 82.880 26.380 83.050 28.460 ;
        RECT 83.680 27.960 84.130 28.130 ;
        RECT 83.450 26.750 83.620 27.790 ;
        RECT 84.190 26.750 84.360 27.790 ;
        RECT 84.760 26.380 84.930 28.460 ;
        RECT 82.880 26.210 84.930 26.380 ;
        RECT 85.430 30.720 87.480 30.890 ;
        RECT 85.430 28.640 85.600 30.720 ;
        RECT 86.230 30.210 86.680 30.380 ;
        RECT 86.000 29.000 86.170 30.040 ;
        RECT 86.740 29.000 86.910 30.040 ;
        RECT 87.310 28.640 87.480 30.720 ;
        RECT 85.430 28.460 87.480 28.640 ;
        RECT 85.430 26.380 85.600 28.460 ;
        RECT 86.230 27.960 86.680 28.130 ;
        RECT 86.000 26.750 86.170 27.790 ;
        RECT 86.740 26.750 86.910 27.790 ;
        RECT 87.310 26.380 87.480 28.460 ;
        RECT 85.430 26.210 87.480 26.380 ;
        RECT 87.980 30.720 90.030 30.890 ;
        RECT 87.980 28.640 88.150 30.720 ;
        RECT 88.780 30.210 89.230 30.380 ;
        RECT 88.550 29.000 88.720 30.040 ;
        RECT 89.290 29.000 89.460 30.040 ;
        RECT 89.860 28.640 90.030 30.720 ;
        RECT 87.980 28.460 90.030 28.640 ;
        RECT 87.980 26.380 88.150 28.460 ;
        RECT 88.780 27.960 89.230 28.130 ;
        RECT 88.550 26.750 88.720 27.790 ;
        RECT 89.290 26.750 89.460 27.790 ;
        RECT 89.860 26.380 90.030 28.460 ;
        RECT 87.980 26.210 90.030 26.380 ;
        RECT 90.530 30.720 92.580 30.890 ;
        RECT 90.530 28.640 90.700 30.720 ;
        RECT 91.330 30.210 91.780 30.380 ;
        RECT 91.100 29.000 91.270 30.040 ;
        RECT 91.840 29.000 92.010 30.040 ;
        RECT 92.410 28.640 92.580 30.720 ;
        RECT 90.530 28.460 92.580 28.640 ;
        RECT 90.530 26.380 90.700 28.460 ;
        RECT 91.330 27.960 91.780 28.130 ;
        RECT 91.100 26.750 91.270 27.790 ;
        RECT 91.840 26.750 92.010 27.790 ;
        RECT 92.410 26.380 92.580 28.460 ;
        RECT 90.530 26.210 92.580 26.380 ;
        RECT 93.080 30.720 95.130 30.890 ;
        RECT 93.080 28.640 93.250 30.720 ;
        RECT 93.880 30.210 94.330 30.380 ;
        RECT 93.650 29.000 93.820 30.040 ;
        RECT 94.390 29.000 94.560 30.040 ;
        RECT 94.960 28.640 95.130 30.720 ;
        RECT 93.080 28.460 95.130 28.640 ;
        RECT 93.080 26.380 93.250 28.460 ;
        RECT 93.880 27.960 94.330 28.130 ;
        RECT 93.650 26.750 93.820 27.790 ;
        RECT 94.390 26.750 94.560 27.790 ;
        RECT 94.960 26.380 95.130 28.460 ;
        RECT 93.080 26.210 95.130 26.380 ;
        RECT 95.630 30.720 97.680 30.890 ;
        RECT 95.630 28.640 95.800 30.720 ;
        RECT 96.430 30.210 96.880 30.380 ;
        RECT 96.200 29.000 96.370 30.040 ;
        RECT 96.940 29.000 97.110 30.040 ;
        RECT 97.510 28.640 97.680 30.720 ;
        RECT 95.630 28.460 97.680 28.640 ;
        RECT 95.630 26.380 95.800 28.460 ;
        RECT 96.430 27.960 96.880 28.130 ;
        RECT 96.200 26.750 96.370 27.790 ;
        RECT 96.940 26.750 97.110 27.790 ;
        RECT 97.510 26.380 97.680 28.460 ;
        RECT 95.630 26.210 97.680 26.380 ;
      LAYER met1 ;
        RECT 72.350 42.430 95.660 42.880 ;
        RECT 85.540 42.400 95.660 42.430 ;
        RECT 78.550 41.275 78.950 41.380 ;
        RECT 85.620 41.275 85.910 41.935 ;
        RECT 87.000 41.860 87.290 41.905 ;
        RECT 87.920 41.860 88.210 41.905 ;
        RECT 93.440 41.860 93.730 41.905 ;
        RECT 87.000 41.720 93.730 41.860 ;
        RECT 87.000 41.675 87.290 41.720 ;
        RECT 87.920 41.675 88.210 41.720 ;
        RECT 93.440 41.675 93.730 41.720 ;
        RECT 86.495 41.520 86.785 41.565 ;
        RECT 88.335 41.520 88.625 41.565 ;
        RECT 86.495 41.380 88.625 41.520 ;
        RECT 86.495 41.335 86.785 41.380 ;
        RECT 88.335 41.335 88.625 41.380 ;
        RECT 88.765 41.280 89.155 41.570 ;
        RECT 89.540 41.280 89.975 41.580 ;
        RECT 90.120 41.280 90.510 41.580 ;
        RECT 90.680 41.520 90.970 41.565 ;
        RECT 92.520 41.520 92.810 41.565 ;
        RECT 93.900 41.540 94.190 41.595 ;
        RECT 90.680 41.380 92.810 41.520 ;
        RECT 90.680 41.335 90.970 41.380 ;
        RECT 92.520 41.335 92.810 41.380 ;
        RECT 78.550 41.130 85.910 41.275 ;
        RECT 78.550 41.030 78.950 41.130 ;
        RECT 85.620 40.625 85.910 41.130 ;
        RECT 91.600 41.225 91.890 41.240 ;
        RECT 91.600 40.965 91.940 41.225 ;
        RECT 93.840 41.130 94.250 41.540 ;
        RECT 94.820 41.435 95.110 41.595 ;
        RECT 93.900 40.965 94.190 41.130 ;
        RECT 94.745 41.025 95.155 41.435 ;
        RECT 94.820 40.965 95.110 41.025 ;
        RECT 91.600 40.945 91.890 40.965 ;
        RECT 87.415 40.840 87.705 40.885 ;
        RECT 90.645 40.840 90.935 40.885 ;
        RECT 87.415 40.700 90.935 40.840 ;
        RECT 87.415 40.655 87.705 40.700 ;
        RECT 90.645 40.655 90.935 40.700 ;
        RECT 85.540 40.130 95.660 40.160 ;
        RECT 74.450 39.680 95.660 40.130 ;
        RECT 74.470 38.330 75.080 38.350 ;
        RECT 72.700 37.780 97.950 38.330 ;
        RECT 74.450 37.740 75.080 37.780 ;
        RECT 74.450 36.430 74.900 37.740 ;
        RECT 76.550 37.530 77.350 37.780 ;
        RECT 79.100 37.530 79.900 37.780 ;
        RECT 81.650 37.530 82.450 37.780 ;
        RECT 84.200 37.530 85.000 37.780 ;
        RECT 86.750 37.530 87.550 37.780 ;
        RECT 89.300 37.530 90.100 37.780 ;
        RECT 91.850 37.530 92.650 37.780 ;
        RECT 94.400 37.530 95.200 37.780 ;
        RECT 96.950 37.530 97.750 37.780 ;
        RECT 73.450 34.230 73.750 36.430 ;
        RECT 74.050 34.430 74.900 36.430 ;
        RECT 73.450 33.780 74.050 34.230 ;
        RECT 74.450 33.930 74.900 34.430 ;
        RECT 75.200 35.530 76.000 37.530 ;
        RECT 76.510 35.530 77.350 37.530 ;
        RECT 77.750 35.530 78.550 37.530 ;
        RECT 79.060 35.530 79.900 37.530 ;
        RECT 80.300 35.530 81.100 37.530 ;
        RECT 81.610 35.530 82.450 37.530 ;
        RECT 82.850 35.530 83.650 37.530 ;
        RECT 84.160 35.530 85.000 37.530 ;
        RECT 85.400 35.530 86.200 37.530 ;
        RECT 86.710 35.530 87.550 37.530 ;
        RECT 87.950 35.530 88.750 37.530 ;
        RECT 89.260 35.530 90.100 37.530 ;
        RECT 90.500 35.530 91.300 37.530 ;
        RECT 91.810 35.530 92.650 37.530 ;
        RECT 93.050 35.530 93.850 37.530 ;
        RECT 94.360 35.530 95.200 37.530 ;
        RECT 95.600 35.530 96.400 37.530 ;
        RECT 96.910 35.530 97.750 37.530 ;
        RECT 75.200 34.230 75.600 35.530 ;
        RECT 75.750 34.830 76.750 35.380 ;
        RECT 77.750 34.230 78.150 35.530 ;
        RECT 78.300 34.830 79.300 35.380 ;
        RECT 80.300 34.230 80.700 35.530 ;
        RECT 80.850 34.830 81.850 35.380 ;
        RECT 82.850 34.230 83.250 35.530 ;
        RECT 83.400 34.830 84.400 35.380 ;
        RECT 85.400 34.230 85.800 35.530 ;
        RECT 85.950 34.830 86.950 35.380 ;
        RECT 87.950 34.230 88.350 35.530 ;
        RECT 88.500 34.830 89.500 35.380 ;
        RECT 90.500 34.230 90.900 35.530 ;
        RECT 91.050 34.830 92.050 35.380 ;
        RECT 93.050 34.230 93.450 35.530 ;
        RECT 93.600 34.830 94.600 35.380 ;
        RECT 95.600 34.230 96.000 35.530 ;
        RECT 96.150 34.830 97.150 35.380 ;
        RECT 73.450 32.930 73.750 33.780 ;
        RECT 73.300 32.430 73.900 32.930 ;
        RECT 73.450 28.030 73.750 32.430 ;
        RECT 75.200 32.230 76.000 34.230 ;
        RECT 76.510 32.230 77.300 34.230 ;
        RECT 77.750 32.230 78.550 34.230 ;
        RECT 79.060 32.230 79.850 34.230 ;
        RECT 80.300 32.230 81.100 34.230 ;
        RECT 81.610 32.230 82.400 34.230 ;
        RECT 82.850 32.230 83.650 34.230 ;
        RECT 84.160 32.230 84.950 34.230 ;
        RECT 85.400 32.230 86.200 34.230 ;
        RECT 86.710 32.230 87.500 34.230 ;
        RECT 87.950 32.230 88.750 34.230 ;
        RECT 89.260 32.230 90.050 34.230 ;
        RECT 90.500 32.230 91.300 34.230 ;
        RECT 91.810 32.230 92.600 34.230 ;
        RECT 93.050 32.230 93.850 34.230 ;
        RECT 94.360 32.230 95.150 34.230 ;
        RECT 95.600 32.230 96.400 34.230 ;
        RECT 96.910 32.230 97.700 34.230 ;
        RECT 76.000 31.380 76.500 32.030 ;
        RECT 75.000 30.830 76.500 31.380 ;
        RECT 76.000 30.180 76.500 30.830 ;
        RECT 76.800 31.380 77.300 32.230 ;
        RECT 78.550 31.380 79.050 32.030 ;
        RECT 76.800 30.830 79.050 31.380 ;
        RECT 74.060 29.930 74.290 29.980 ;
        RECT 74.550 29.930 74.900 30.130 ;
        RECT 76.800 30.030 77.300 30.830 ;
        RECT 78.550 30.180 79.050 30.830 ;
        RECT 79.350 31.380 79.850 32.230 ;
        RECT 81.100 31.380 81.600 32.030 ;
        RECT 81.900 31.380 82.400 32.230 ;
        RECT 83.650 31.380 84.150 32.030 ;
        RECT 79.350 30.830 81.600 31.380 ;
        RECT 81.850 30.830 84.150 31.380 ;
        RECT 79.350 30.030 79.850 30.830 ;
        RECT 81.100 30.180 81.600 30.830 ;
        RECT 81.900 30.030 82.400 30.830 ;
        RECT 83.650 30.180 84.150 30.830 ;
        RECT 84.450 31.380 84.950 32.230 ;
        RECT 86.200 31.380 86.700 32.030 ;
        RECT 87.000 31.380 87.500 32.230 ;
        RECT 88.750 31.380 89.250 32.030 ;
        RECT 84.450 30.830 86.700 31.380 ;
        RECT 86.950 30.830 89.250 31.380 ;
        RECT 84.450 30.030 84.950 30.830 ;
        RECT 86.200 30.180 86.700 30.830 ;
        RECT 87.000 30.030 87.500 30.830 ;
        RECT 88.750 30.180 89.250 30.830 ;
        RECT 89.550 31.380 90.050 32.230 ;
        RECT 91.300 31.380 91.800 32.030 ;
        RECT 92.100 31.380 92.600 32.230 ;
        RECT 93.850 31.380 94.350 32.030 ;
        RECT 89.550 30.830 91.800 31.380 ;
        RECT 92.050 30.830 94.350 31.380 ;
        RECT 89.550 30.030 90.050 30.830 ;
        RECT 91.300 30.180 91.800 30.830 ;
        RECT 92.100 30.030 92.600 30.830 ;
        RECT 93.850 30.180 94.350 30.830 ;
        RECT 94.650 31.380 95.150 32.230 ;
        RECT 96.400 31.380 96.900 32.030 ;
        RECT 97.200 31.380 97.700 32.230 ;
        RECT 94.650 30.830 96.900 31.380 ;
        RECT 97.150 30.830 98.000 31.380 ;
        RECT 94.650 30.030 95.150 30.830 ;
        RECT 96.400 30.180 96.900 30.830 ;
        RECT 97.200 30.030 97.700 30.830 ;
        RECT 74.050 28.030 74.900 29.930 ;
        RECT 73.470 27.980 73.700 28.030 ;
        RECT 74.060 27.980 74.290 28.030 ;
        RECT 73.600 27.380 74.150 27.830 ;
        RECT 72.370 26.580 72.980 26.610 ;
        RECT 74.550 26.580 74.900 28.030 ;
        RECT 75.200 30.020 75.950 30.030 ;
        RECT 76.550 30.020 77.300 30.030 ;
        RECT 75.200 29.030 76.000 30.020 ;
        RECT 75.200 27.780 75.600 29.030 ;
        RECT 75.770 29.020 76.000 29.030 ;
        RECT 76.510 29.030 77.300 30.020 ;
        RECT 77.750 30.020 78.500 30.030 ;
        RECT 79.100 30.020 79.850 30.030 ;
        RECT 77.750 29.030 78.550 30.020 ;
        RECT 76.510 29.020 76.740 29.030 ;
        RECT 75.750 27.930 76.750 28.480 ;
        RECT 77.050 27.780 77.350 28.030 ;
        RECT 75.200 27.770 75.950 27.780 ;
        RECT 76.550 27.770 77.350 27.780 ;
        RECT 75.200 26.780 76.000 27.770 ;
        RECT 75.770 26.770 76.000 26.780 ;
        RECT 76.510 26.770 77.350 27.770 ;
        RECT 77.750 27.780 78.150 29.030 ;
        RECT 78.320 29.020 78.550 29.030 ;
        RECT 79.060 29.030 79.850 30.020 ;
        RECT 80.300 30.020 81.050 30.030 ;
        RECT 81.650 30.020 82.400 30.030 ;
        RECT 80.300 29.030 81.100 30.020 ;
        RECT 79.060 29.020 79.290 29.030 ;
        RECT 78.300 27.930 79.300 28.480 ;
        RECT 79.600 27.780 79.900 28.030 ;
        RECT 77.750 27.770 78.500 27.780 ;
        RECT 79.100 27.770 79.900 27.780 ;
        RECT 77.750 26.780 78.550 27.770 ;
        RECT 78.320 26.770 78.550 26.780 ;
        RECT 79.060 26.770 79.900 27.770 ;
        RECT 80.300 27.780 80.700 29.030 ;
        RECT 80.870 29.020 81.100 29.030 ;
        RECT 81.610 29.030 82.400 30.020 ;
        RECT 82.850 30.020 83.600 30.030 ;
        RECT 84.200 30.020 84.950 30.030 ;
        RECT 82.850 29.030 83.650 30.020 ;
        RECT 81.610 29.020 81.840 29.030 ;
        RECT 80.850 27.930 81.850 28.480 ;
        RECT 82.150 27.780 82.450 28.030 ;
        RECT 80.300 27.770 81.050 27.780 ;
        RECT 81.650 27.770 82.450 27.780 ;
        RECT 80.300 26.780 81.100 27.770 ;
        RECT 80.870 26.770 81.100 26.780 ;
        RECT 81.610 26.770 82.450 27.770 ;
        RECT 82.850 27.780 83.250 29.030 ;
        RECT 83.420 29.020 83.650 29.030 ;
        RECT 84.160 29.030 84.950 30.020 ;
        RECT 85.400 30.020 86.150 30.030 ;
        RECT 86.750 30.020 87.500 30.030 ;
        RECT 85.400 29.030 86.200 30.020 ;
        RECT 84.160 29.020 84.390 29.030 ;
        RECT 83.400 27.930 84.400 28.480 ;
        RECT 84.700 27.780 85.000 28.030 ;
        RECT 82.850 27.770 83.600 27.780 ;
        RECT 84.200 27.770 85.000 27.780 ;
        RECT 82.850 26.780 83.650 27.770 ;
        RECT 83.420 26.770 83.650 26.780 ;
        RECT 84.160 26.770 85.000 27.770 ;
        RECT 85.400 27.780 85.800 29.030 ;
        RECT 85.970 29.020 86.200 29.030 ;
        RECT 86.710 29.030 87.500 30.020 ;
        RECT 87.950 30.020 88.700 30.030 ;
        RECT 89.300 30.020 90.050 30.030 ;
        RECT 87.950 29.030 88.750 30.020 ;
        RECT 86.710 29.020 86.940 29.030 ;
        RECT 85.950 27.930 86.950 28.480 ;
        RECT 87.250 27.780 87.550 28.030 ;
        RECT 85.400 27.770 86.150 27.780 ;
        RECT 86.750 27.770 87.550 27.780 ;
        RECT 85.400 26.780 86.200 27.770 ;
        RECT 85.970 26.770 86.200 26.780 ;
        RECT 86.710 26.770 87.550 27.770 ;
        RECT 87.950 27.780 88.350 29.030 ;
        RECT 88.520 29.020 88.750 29.030 ;
        RECT 89.260 29.030 90.050 30.020 ;
        RECT 90.500 30.020 91.250 30.030 ;
        RECT 91.850 30.020 92.600 30.030 ;
        RECT 90.500 29.030 91.300 30.020 ;
        RECT 89.260 29.020 89.490 29.030 ;
        RECT 88.500 27.930 89.500 28.480 ;
        RECT 89.800 27.780 90.100 28.030 ;
        RECT 87.950 27.770 88.700 27.780 ;
        RECT 89.300 27.770 90.100 27.780 ;
        RECT 87.950 26.780 88.750 27.770 ;
        RECT 88.520 26.770 88.750 26.780 ;
        RECT 89.260 26.770 90.100 27.770 ;
        RECT 90.500 27.780 90.900 29.030 ;
        RECT 91.070 29.020 91.300 29.030 ;
        RECT 91.810 29.030 92.600 30.020 ;
        RECT 93.050 30.020 93.800 30.030 ;
        RECT 94.400 30.020 95.150 30.030 ;
        RECT 93.050 29.030 93.850 30.020 ;
        RECT 91.810 29.020 92.040 29.030 ;
        RECT 91.050 27.930 92.050 28.480 ;
        RECT 92.350 27.780 92.650 28.030 ;
        RECT 90.500 27.770 91.250 27.780 ;
        RECT 91.850 27.770 92.650 27.780 ;
        RECT 90.500 26.780 91.300 27.770 ;
        RECT 91.070 26.770 91.300 26.780 ;
        RECT 91.810 26.770 92.650 27.770 ;
        RECT 93.050 27.780 93.450 29.030 ;
        RECT 93.620 29.020 93.850 29.030 ;
        RECT 94.360 29.030 95.150 30.020 ;
        RECT 95.600 30.020 96.350 30.030 ;
        RECT 96.950 30.020 97.700 30.030 ;
        RECT 95.600 29.030 96.400 30.020 ;
        RECT 94.360 29.020 94.590 29.030 ;
        RECT 93.600 27.930 94.600 28.480 ;
        RECT 94.900 27.780 95.200 28.030 ;
        RECT 93.050 27.770 93.800 27.780 ;
        RECT 94.400 27.770 95.200 27.780 ;
        RECT 93.050 26.780 93.850 27.770 ;
        RECT 93.620 26.770 93.850 26.780 ;
        RECT 94.360 26.770 95.200 27.770 ;
        RECT 95.600 27.780 96.000 29.030 ;
        RECT 96.170 29.020 96.400 29.030 ;
        RECT 96.910 29.030 97.700 30.020 ;
        RECT 96.910 29.020 97.140 29.030 ;
        RECT 96.150 27.930 97.150 28.480 ;
        RECT 97.450 27.780 97.750 28.030 ;
        RECT 95.600 27.770 96.350 27.780 ;
        RECT 96.950 27.770 97.750 27.780 ;
        RECT 95.600 26.780 96.400 27.770 ;
        RECT 96.170 26.770 96.400 26.780 ;
        RECT 96.910 26.770 97.750 27.770 ;
        RECT 76.550 26.580 77.350 26.770 ;
        RECT 79.100 26.580 79.900 26.770 ;
        RECT 81.650 26.580 82.450 26.770 ;
        RECT 84.200 26.580 85.000 26.770 ;
        RECT 86.750 26.580 87.550 26.770 ;
        RECT 89.300 26.580 90.100 26.770 ;
        RECT 91.850 26.580 92.650 26.770 ;
        RECT 94.400 26.580 95.200 26.770 ;
        RECT 96.950 26.580 97.750 26.770 ;
        RECT 72.370 26.030 97.950 26.580 ;
        RECT 72.370 26.000 72.980 26.030 ;
      LAYER met2 ;
        RECT 72.400 42.380 72.950 42.930 ;
        RECT 80.480 42.435 81.070 43.025 ;
        RECT 78.600 40.980 78.900 41.430 ;
        RECT 74.500 39.630 75.050 40.180 ;
        RECT 80.655 38.535 80.900 42.435 ;
        RECT 82.480 42.340 83.070 42.840 ;
        RECT 82.650 41.565 82.905 42.340 ;
        RECT 88.815 41.565 89.105 41.620 ;
        RECT 82.650 41.310 89.105 41.565 ;
        RECT 88.815 41.230 89.105 41.310 ;
        RECT 89.590 41.230 89.880 41.630 ;
        RECT 90.170 41.230 90.460 41.630 ;
        RECT 89.605 39.045 89.850 41.230 ;
        RECT 90.195 39.810 90.430 41.230 ;
        RECT 91.650 40.935 91.910 41.255 ;
        RECT 93.840 41.130 94.250 41.540 ;
        RECT 94.745 41.025 95.155 41.435 ;
        RECT 90.160 39.420 90.460 39.810 ;
        RECT 89.530 38.745 89.920 39.045 ;
        RECT 91.655 38.535 91.900 40.935 ;
        RECT 74.470 37.740 75.080 38.350 ;
        RECT 80.655 38.290 91.900 38.535 ;
        RECT 73.350 34.830 97.950 35.380 ;
        RECT 73.350 32.380 73.850 34.830 ;
        RECT 74.355 33.125 74.855 33.145 ;
        RECT 74.330 28.380 74.880 33.125 ;
        RECT 75.200 30.780 75.950 31.430 ;
        RECT 81.900 30.780 82.650 31.430 ;
        RECT 87.000 30.780 87.750 31.430 ;
        RECT 92.100 30.780 92.850 31.430 ;
        RECT 97.200 30.780 97.950 31.430 ;
        RECT 75.750 28.380 97.950 28.480 ;
        RECT 72.700 28.030 97.950 28.380 ;
        RECT 73.650 27.330 74.100 28.030 ;
        RECT 75.750 27.930 97.950 28.030 ;
        RECT 72.370 26.000 72.980 26.610 ;
      LAYER met3 ;
        RECT 142.360 133.650 142.740 133.660 ;
        RECT 147.470 133.650 147.850 133.690 ;
        RECT 142.360 133.350 147.850 133.650 ;
        RECT 142.360 133.340 142.740 133.350 ;
        RECT 147.470 133.310 147.850 133.350 ;
        RECT 0.950 46.060 2.550 46.300 ;
        RECT 0.950 44.945 75.305 46.060 ;
        RECT 0.950 44.700 2.550 44.945 ;
        RECT 49.005 43.155 50.495 43.425 ;
        RECT 72.400 43.155 72.950 43.180 ;
        RECT 49.005 42.905 72.955 43.155 ;
        RECT 49.005 42.405 73.000 42.905 ;
        RECT 49.005 42.145 72.955 42.405 ;
        RECT 74.190 42.145 75.305 44.945 ;
        RECT 76.510 45.935 157.230 45.940 ;
        RECT 76.510 45.260 157.255 45.935 ;
        RECT 76.510 45.255 157.230 45.260 ;
        RECT 49.005 41.875 50.495 42.145 ;
        RECT 72.400 26.030 72.950 42.145 ;
        RECT 74.500 40.155 75.050 42.145 ;
        RECT 76.510 42.060 77.195 45.255 ;
        RECT 78.500 43.050 79.050 43.180 ;
        RECT 80.500 43.050 81.050 43.180 ;
        RECT 82.500 43.050 83.050 43.180 ;
        RECT 78.400 42.400 79.150 43.050 ;
        RECT 80.400 42.400 81.150 43.050 ;
        RECT 82.400 42.400 83.150 43.050 ;
        RECT 78.500 42.180 79.050 42.400 ;
        RECT 80.500 42.180 81.050 42.400 ;
        RECT 82.500 42.180 83.050 42.400 ;
        RECT 92.350 42.205 95.125 42.555 ;
        RECT 74.450 39.655 75.100 40.155 ;
        RECT 74.500 37.770 75.050 39.655 ;
        RECT 76.550 33.125 77.100 42.060 ;
        RECT 78.595 41.405 78.920 42.180 ;
        RECT 78.550 41.005 78.950 41.405 ;
        RECT 74.330 32.575 77.100 33.125 ;
        RECT 75.150 31.300 76.000 31.405 ;
        RECT 78.595 31.300 78.920 41.005 ;
        RECT 82.100 39.440 90.485 39.790 ;
        RECT 82.100 31.405 82.450 39.440 ;
        RECT 87.200 38.720 89.900 39.070 ;
        RECT 87.200 31.405 87.550 38.720 ;
        RECT 92.350 31.405 92.700 42.205 ;
        RECT 93.870 39.200 94.220 41.510 ;
        RECT 94.775 41.055 95.125 42.205 ;
        RECT 93.870 38.850 97.800 39.200 ;
        RECT 97.450 31.405 97.800 38.850 ;
        RECT 75.150 30.975 78.920 31.300 ;
        RECT 75.150 30.805 76.000 30.975 ;
        RECT 81.850 30.805 82.700 31.405 ;
        RECT 86.950 30.805 87.800 31.405 ;
        RECT 92.050 30.805 92.900 31.405 ;
        RECT 97.150 30.805 98.000 31.405 ;
      LAYER met4 ;
        RECT 3.990 222.300 4.290 224.760 ;
        RECT 7.670 224.000 7.970 224.760 ;
        RECT 11.350 224.000 11.650 224.760 ;
        RECT 15.030 224.000 15.330 224.760 ;
        RECT 18.710 224.000 19.010 224.760 ;
        RECT 22.390 224.000 22.690 224.760 ;
        RECT 26.070 224.000 26.370 224.760 ;
        RECT 29.750 224.000 30.050 224.760 ;
        RECT 33.430 224.000 33.730 224.760 ;
        RECT 37.110 224.000 37.410 224.760 ;
        RECT 40.790 224.000 41.090 224.760 ;
        RECT 44.470 224.000 44.770 224.760 ;
        RECT 48.150 224.000 48.450 224.760 ;
        RECT 51.830 224.000 52.130 224.760 ;
        RECT 55.510 224.000 55.810 224.760 ;
        RECT 59.190 224.000 59.490 224.760 ;
        RECT 62.870 224.000 63.170 224.760 ;
        RECT 66.550 224.000 66.850 224.760 ;
        RECT 70.230 224.000 70.530 224.760 ;
        RECT 73.910 224.000 74.210 224.760 ;
        RECT 77.590 224.000 77.890 224.760 ;
        RECT 81.270 224.000 81.570 224.760 ;
        RECT 84.950 224.000 85.250 224.760 ;
        RECT 6.100 222.300 86.350 224.000 ;
        RECT 3.990 222.000 86.350 222.300 ;
        RECT 1.000 27.155 2.500 220.760 ;
        RECT 6.100 220.550 86.350 222.000 ;
        RECT 0.995 25.700 2.505 27.155 ;
        RECT 0.995 25.695 1.000 25.700 ;
        RECT 2.500 25.695 2.505 25.700 ;
        RECT 49.000 14.755 50.500 220.550 ;
        RECT 88.630 68.250 88.930 224.760 ;
        RECT 142.385 133.335 142.715 133.665 ;
        RECT 78.600 67.950 88.930 68.250 ;
        RECT 78.600 44.200 78.900 67.950 ;
        RECT 142.400 52.000 142.700 133.335 ;
        RECT 80.550 51.700 142.700 52.000 ;
        RECT 80.550 44.200 80.850 51.700 ;
        RECT 143.830 50.200 144.130 224.760 ;
        RECT 147.510 133.665 147.810 224.760 ;
        RECT 147.495 133.335 147.825 133.665 ;
        RECT 82.550 49.900 144.130 50.200 ;
        RECT 82.550 44.200 82.850 49.900 ;
        RECT 143.830 49.800 144.130 49.900 ;
        RECT 78.450 43.055 79.100 44.200 ;
        RECT 80.450 43.055 81.100 44.200 ;
        RECT 82.450 43.055 83.100 44.200 ;
        RECT 78.445 42.395 79.105 43.055 ;
        RECT 80.445 42.395 81.105 43.055 ;
        RECT 82.445 42.395 83.105 43.055 ;
        RECT 78.450 42.375 79.100 42.395 ;
        RECT 48.995 13.300 50.505 14.755 ;
        RECT 48.995 13.295 49.000 13.300 ;
        RECT 50.500 13.295 50.505 13.300 ;
        RECT 156.545 1.000 157.230 45.940 ;
  END
END tt_um_obriensp_pll
END LIBRARY

