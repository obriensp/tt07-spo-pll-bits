magic
tech sky130A
magscale 1 2
timestamp 1717213418
<< metal1 >>
rect 0 -770 200 -570
rect 1530 -720 1870 -570
rect 3400 -890 3600 -870
rect 10 -1050 20 -890
rect 180 -1050 190 -890
rect 3400 -1050 3420 -890
rect 3580 -1050 3600 -890
rect 3400 -1070 3600 -1050
rect 0 -1380 200 -1180
rect 1800 -1380 2000 -1180
rect 3400 -1540 3600 -1520
rect 10 -1700 20 -1540
rect 180 -1700 190 -1540
rect 3400 -1700 3420 -1540
rect 3580 -1700 3600 -1540
rect 3400 -1720 3600 -1700
rect 0 -2000 200 -1800
rect 1520 -2000 1860 -1910
<< via1 >>
rect 20 -1050 180 -890
rect 3420 -1050 3580 -890
rect 20 -1700 180 -1540
rect 3420 -1700 3580 -1540
<< metal2 >>
rect 20 -890 180 -880
rect 3420 -890 3580 -880
rect 1630 -935 1710 -930
rect 1626 -1005 1635 -935
rect 1705 -1005 1714 -935
rect 20 -1060 180 -1050
rect 20 -1540 180 -1530
rect 1630 -1580 1710 -1005
rect 3420 -1060 3580 -1050
rect 1630 -1669 1710 -1660
rect 3420 -1540 3580 -1530
rect 20 -1710 180 -1700
rect 3420 -1710 3580 -1700
<< via2 >>
rect 20 -1050 180 -890
rect 1635 -1005 1705 -935
rect 20 -1700 180 -1540
rect 3420 -1050 3580 -890
rect 1630 -1660 1710 -1580
rect 3420 -1700 3580 -1540
<< metal3 >>
rect 10 -890 190 -885
rect 10 -1050 20 -890
rect 180 -930 190 -890
rect 3410 -890 3590 -885
rect 3410 -930 3420 -890
rect 180 -1010 1480 -930
rect 1630 -935 3420 -930
rect 1630 -1005 1635 -935
rect 1705 -1005 3420 -935
rect 1630 -1010 3420 -1005
rect 180 -1050 190 -1010
rect 10 -1055 190 -1050
rect 1400 -1430 1480 -1010
rect 3410 -1050 3420 -1010
rect 3580 -1050 3590 -890
rect 3410 -1055 3590 -1050
rect 1400 -1510 3270 -1430
rect 10 -1540 190 -1535
rect 10 -1700 20 -1540
rect 180 -1580 190 -1540
rect 1625 -1580 1715 -1575
rect 180 -1660 1630 -1580
rect 1710 -1660 1715 -1580
rect 3190 -1580 3270 -1510
rect 3410 -1540 3590 -1535
rect 3410 -1580 3420 -1540
rect 3190 -1660 3420 -1580
rect 180 -1700 190 -1660
rect 1625 -1665 1715 -1660
rect 10 -1705 190 -1700
rect 3410 -1700 3420 -1660
rect 3580 -1700 3590 -1540
rect 3410 -1705 3590 -1700
use latch  x2
timestamp 1717213418
transform 1 0 -1040 0 1 650
box 1040 -2650 2840 -1220
use latch  x3
timestamp 1717213418
transform 1 0 760 0 1 650
box 1040 -2650 2840 -1220
<< labels >>
flabel metal1 3400 -1070 3600 -870 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 3400 -1720 3600 -1520 0 FreeSans 256 0 0 0 out_n
port 3 nsew
flabel metal1 0 -1380 200 -1180 0 FreeSans 256 0 0 0 clk
port 5 nsew
flabel metal1 0 -770 200 -570 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 1800 -1380 2000 -1180 0 FreeSans 256 0 0 0 clk_n
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vss
port 1 nsew
<< end >>
