magic
tech sky130A
magscale 1 2
timestamp 1717079806
<< error_s >>
rect 5160 3780 5546 3860
rect 4930 1776 4988 1782
rect 5078 1776 5136 1782
rect 4782 1146 5292 1776
rect 5004 1144 5062 1146
rect 4930 -54 4988 -48
rect 5078 -54 5136 -48
rect 4782 -684 5292 -54
rect 5004 -686 5062 -684
rect 4800 -2240 5292 -1818
rect 4822 -2364 4828 -2342
rect 4942 -2354 4976 -2240
rect 5090 -2354 5124 -2240
rect 5204 -2340 5238 -2240
rect 4794 -2392 4800 -2370
<< viali >>
rect 5292 4478 5450 4512
rect 5196 3913 5230 4415
rect 5722 4268 5880 4302
rect 5942 3912 5976 4206
rect 5292 3816 5450 3850
rect 5722 3816 5880 3850
rect 4932 -2204 5506 -2170
rect 5782 -2204 6076 -2170
<< metal1 >>
rect 5480 4580 5680 4780
rect 5178 4512 5464 4524
rect 5178 4478 5292 4512
rect 5450 4478 5464 4512
rect 5178 4466 5464 4478
rect 5178 4415 5296 4466
rect 5178 4274 5196 4415
rect 4484 4074 4490 4274
rect 4690 4074 5196 4274
rect 5178 3913 5196 4074
rect 5230 4402 5296 4415
rect 5230 4000 5350 4402
rect 5550 4260 5620 4580
rect 5400 4214 5620 4260
rect 5694 4302 5996 4324
rect 5694 4268 5722 4302
rect 5880 4268 5996 4302
rect 5694 4252 5996 4268
rect 5230 3913 5296 4000
rect 5400 3990 5780 4214
rect 5890 4206 5996 4252
rect 5890 4190 5942 4206
rect 5822 3992 5942 4190
rect 5848 3990 5942 3992
rect 5178 3862 5296 3913
rect 5330 3890 5840 3960
rect 5890 3912 5942 3990
rect 5976 4148 5996 4206
rect 5976 3948 6520 4148
rect 6720 3948 6726 4148
rect 5976 3912 5996 3948
rect 5178 3850 5460 3862
rect 5178 3816 5292 3850
rect 5450 3816 5460 3850
rect 5178 3804 5460 3816
rect 5550 3736 5620 3890
rect 5890 3860 5996 3912
rect 5694 3850 5996 3860
rect 5694 3816 5722 3850
rect 5880 3816 5996 3850
rect 5694 3806 5996 3816
rect 5694 3796 5994 3806
rect 5148 3536 5158 3736
rect 5358 3536 5368 3736
rect 5474 3536 5484 3736
rect 5684 3536 5694 3736
rect 5788 3536 5798 3736
rect 5998 3536 6008 3736
rect 4494 2420 4504 2624
rect 4728 2420 4738 2624
rect 4120 1912 4130 2112
rect 4330 1912 4340 2112
rect 4792 1914 4802 2114
rect 5002 1914 5012 2114
rect 5148 1706 5158 1906
rect 5358 1706 5368 1906
rect 5480 1700 5690 2110
rect 6110 1912 6120 2112
rect 6320 1912 6330 2112
rect 6508 1912 6518 2112
rect 6718 1912 6728 2112
rect 5788 1706 5798 1906
rect 5998 1706 6008 1906
rect 4494 590 4504 794
rect 4728 590 4738 794
rect 4120 82 4130 282
rect 4330 82 4340 282
rect 4792 84 4802 284
rect 5002 84 5012 284
rect 5148 -124 5158 76
rect 5358 -124 5368 76
rect 5480 -130 5690 280
rect 6110 82 6120 282
rect 6320 82 6330 282
rect 6508 82 6518 282
rect 6718 82 6728 282
rect 5788 -124 5798 76
rect 5998 -124 6008 76
rect 4494 -1240 4504 -1036
rect 4728 -1240 4738 -1036
rect 4120 -1748 4130 -1548
rect 4330 -1748 4340 -1548
rect 4792 -1746 4802 -1546
rect 5002 -1746 5012 -1546
rect 4900 -1900 5010 -1746
rect 5476 -1750 5486 -1550
rect 5686 -1750 5696 -1550
rect 6110 -1748 6120 -1548
rect 6320 -1748 6330 -1548
rect 6508 -1748 6518 -1548
rect 6718 -1748 6728 -1548
rect 4900 -2000 6000 -1900
rect 6190 -1980 6280 -1748
rect 4490 -2060 4690 -2054
rect 4120 -2200 4320 -2194
rect 4120 -2880 4320 -2400
rect 4900 -2070 4990 -2000
rect 5020 -2160 5410 -2060
rect 5450 -2070 5540 -2000
rect 5800 -2150 5990 -2050
rect 6030 -2070 6280 -1980
rect 4690 -2170 5520 -2160
rect 4690 -2204 4932 -2170
rect 5506 -2204 5520 -2170
rect 4690 -2220 5520 -2204
rect 5680 -2170 6720 -2150
rect 5680 -2204 5782 -2170
rect 6076 -2204 6720 -2170
rect 5680 -2210 6720 -2204
rect 5680 -2220 6520 -2210
rect 4490 -2370 4690 -2260
rect 4490 -2570 4800 -2370
rect 4600 -2880 4800 -2570
rect 5090 -2450 5290 -2444
rect 5090 -2880 5290 -2650
rect 5530 -2460 5730 -2454
rect 5530 -2880 5730 -2660
rect 6010 -2690 6140 -2490
rect 6340 -2690 6346 -2490
rect 6010 -2880 6210 -2690
rect 6520 -2880 6720 -2410
<< via1 >>
rect 4490 4074 4690 4274
rect 6520 3948 6720 4148
rect 5158 3536 5358 3736
rect 5484 3536 5684 3736
rect 5798 3536 5998 3736
rect 4504 2420 4728 2624
rect 4130 1912 4330 2112
rect 4802 1914 5002 2114
rect 5158 1706 5358 1906
rect 6120 1912 6320 2112
rect 6518 1912 6718 2112
rect 5798 1706 5998 1906
rect 4504 590 4728 794
rect 4130 82 4330 282
rect 4802 84 5002 284
rect 5158 -124 5358 76
rect 6120 82 6320 282
rect 6518 82 6718 282
rect 5798 -124 5998 76
rect 4504 -1240 4728 -1036
rect 4130 -1748 4330 -1548
rect 4802 -1746 5002 -1546
rect 5486 -1750 5686 -1550
rect 6120 -1748 6320 -1548
rect 6518 -1748 6718 -1548
rect 4120 -2400 4320 -2200
rect 4490 -2260 4690 -2060
rect 6520 -2410 6720 -2210
rect 5090 -2650 5290 -2450
rect 5530 -2660 5730 -2460
rect 6140 -2690 6340 -2490
<< metal2 >>
rect 4490 4274 4690 4280
rect 4490 2634 4690 4074
rect 6520 4148 6720 4154
rect 5780 3746 5980 3750
rect 5158 3740 5358 3746
rect 5090 3736 5358 3740
rect 5090 3536 5158 3736
rect 5090 3526 5358 3536
rect 5484 3736 5684 3746
rect 5484 3526 5684 3536
rect 5780 3736 5998 3746
rect 5780 3536 5798 3736
rect 5780 3526 5998 3536
rect 4490 2624 4728 2634
rect 4120 2122 4320 2520
rect 4490 2420 4504 2624
rect 4490 2410 4728 2420
rect 4120 2112 4330 2122
rect 4120 1912 4130 2112
rect 4120 1902 4330 1912
rect 4120 292 4320 1902
rect 4490 804 4690 2410
rect 4802 2114 5002 2124
rect 4490 794 4728 804
rect 4490 590 4504 794
rect 4490 580 4728 590
rect 4120 282 4330 292
rect 4120 82 4130 282
rect 4120 72 4330 82
rect 4120 -1538 4320 72
rect 4490 -1026 4690 580
rect 4802 284 5002 1914
rect 4490 -1036 4728 -1026
rect 4490 -1240 4504 -1036
rect 4490 -1250 4728 -1240
rect 4120 -1548 4330 -1538
rect 4120 -1748 4130 -1548
rect 4120 -1758 4330 -1748
rect 4120 -2200 4320 -1758
rect 4490 -2060 4690 -1250
rect 4802 -1546 5002 84
rect 4802 -1756 5002 -1746
rect 5090 1916 5290 3526
rect 5780 1916 5980 3526
rect 6120 2112 6320 2124
rect 6520 2122 6720 3948
rect 5090 1906 5358 1916
rect 5090 1706 5158 1906
rect 5090 1696 5358 1706
rect 5780 1906 5998 1916
rect 5780 1706 5798 1906
rect 5780 1696 5998 1706
rect 5090 86 5290 1696
rect 5780 86 5980 1696
rect 6120 282 6320 1912
rect 6518 2112 6720 2122
rect 6718 1912 6720 2112
rect 6518 1902 6720 1912
rect 6520 292 6720 1902
rect 5090 76 5358 86
rect 5090 -124 5158 76
rect 5090 -134 5358 -124
rect 5780 76 5998 86
rect 5780 -124 5798 76
rect 5780 -134 5998 -124
rect 4114 -2400 4120 -2200
rect 4320 -2400 4326 -2200
rect 4484 -2260 4490 -2060
rect 4690 -2260 4696 -2060
rect 5090 -2450 5290 -134
rect 5486 -1550 5686 -1540
rect 5486 -1760 5686 -1750
rect 5780 -2330 5980 -134
rect 6120 -1540 6320 82
rect 6518 282 6720 292
rect 6718 82 6720 282
rect 6518 72 6720 82
rect 6520 -1538 6720 72
rect 6120 -1548 6340 -1540
rect 6320 -1748 6340 -1548
rect 6120 -1758 6340 -1748
rect 6518 -1548 6720 -1538
rect 6718 -1748 6720 -1548
rect 6518 -1758 6720 -1748
rect 5084 -2650 5090 -2450
rect 5290 -2650 5296 -2450
rect 5530 -2460 5980 -2330
rect 5524 -2660 5530 -2460
rect 5730 -2530 5980 -2460
rect 6140 -2490 6340 -1758
rect 6520 -2210 6720 -1758
rect 6514 -2410 6520 -2210
rect 6720 -2410 6726 -2210
rect 5730 -2660 5736 -2530
rect 6140 -2696 6340 -2690
<< via2 >>
rect 5484 3536 5684 3736
rect 5486 -1750 5686 -1550
<< metal3 >>
rect 5474 3736 5694 3741
rect 5474 3536 5484 3736
rect 5684 3536 5694 3736
rect 5474 3531 5694 3536
rect 5548 -1545 5612 3531
rect 5476 -1550 5696 -1545
rect 5476 -1750 5486 -1550
rect 5686 -1750 5696 -1550
rect 5476 -1755 5696 -1750
rect 5548 -1760 5612 -1755
use sky130_fd_pr__nfet_01v8_64QSBY  sky130_fd_pr__nfet_01v8_64QSBY_0
timestamp 1716528727
transform 1 0 5801 0 1 4059
box -211 -279 211 279
use delay_stage  x1
timestamp 1717029282
transform 1 0 3672 0 1 156
box 1110 -2670 1620 -210
use delay_stage  x2
timestamp 1717029282
transform 1 0 3672 0 1 1986
box 1110 -2670 1620 -210
use delay_stage  x3
timestamp 1717029282
transform 1 0 3672 0 1 3816
box 1110 -2670 1620 -210
use sky130_fd_pr__pfet_01v8_LGAKDL  XM2
timestamp 1717042859
transform 1 0 5371 0 1 4164
box -211 -384 211 384
use sky130_fd_pr__pfet_01v8_XGAKDL  XM5
timestamp 1716531588
transform 0 1 5219 -1 0 -2029
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_64QSBY  XM6
timestamp 1716528727
transform 0 -1 5929 1 0 -2029
box -211 -279 211 279
<< labels >>
flabel metal1 5480 4580 5680 4780 0 FreeSans 256 0 0 0 out
port 5 nsew
flabel metal1 4120 -2880 4320 -2680 0 FreeSans 256 0 0 0 vss
flabel metal1 6520 -2880 6720 -2680 0 FreeSans 256 0 0 0 vss
port 6 nsew
flabel metal1 5090 -2880 5290 -2680 0 FreeSans 256 0 0 0 s0
port 3 nsew
flabel metal1 4600 -2880 4800 -2680 0 FreeSans 256 0 0 0 vdd
port 1 nsew
flabel metal1 5530 -2880 5730 -2680 0 FreeSans 256 0 0 0 s1
port 4 nsew
flabel metal1 6010 -2880 6210 -2680 0 FreeSans 256 0 0 0 vcont
port 2 nsew
flabel metal1 5480 -130 5690 280 0 FreeSans 160 0 0 0 stage_0_out
flabel metal1 5480 1700 5690 2110 0 FreeSans 160 0 0 0 stage_1_out
<< end >>
