magic
tech sky130A
magscale 1 2
timestamp 1717195371
<< metal1 >>
rect 23470 13280 23790 13290
rect 23470 12980 23480 13280
rect 23780 12980 25840 13280
rect 23470 12970 23790 12980
rect 25570 12640 25680 12980
rect 19962 10490 20162 10496
rect 19562 8810 19762 8816
rect 19562 7516 19762 8610
rect 19962 7516 20162 10290
rect 23520 8860 23840 8870
rect 23520 8560 23530 8860
rect 23830 8560 25120 8860
rect 23520 8550 23840 8560
rect 25690 7720 25910 7730
rect 25690 7540 25710 7720
rect 25890 7540 25910 7720
rect 25690 7510 25910 7540
<< via1 >>
rect 23480 12980 23780 13280
rect 19962 10290 20162 10490
rect 19562 8610 19762 8810
rect 23530 8560 23830 8860
rect 21700 7540 21820 7660
rect 23070 7570 23190 7690
rect 25710 7540 25890 7720
<< metal2 >>
rect 25360 17168 25440 17180
rect 25360 17112 25372 17168
rect 25428 17112 25440 17168
rect 25360 17100 25440 17112
rect 25370 14500 25430 17100
rect 25920 16368 26000 16380
rect 25920 16312 25932 16368
rect 25988 16312 26000 16368
rect 25920 16300 26000 16312
rect 25930 14530 25990 16300
rect 25930 14461 25990 14470
rect 25370 14431 25430 14440
rect 23470 13280 23790 13290
rect 23470 12980 23480 13280
rect 23780 12980 23790 13280
rect 23470 12970 23790 12980
rect 23480 10550 23780 12970
rect 23470 10535 23790 10550
rect 19950 10490 20170 10500
rect 19950 10290 19962 10490
rect 20162 10290 20170 10490
rect 19950 10280 20170 10290
rect 23470 10245 23485 10535
rect 23775 10245 23790 10535
rect 23470 10230 23790 10245
rect 23520 8860 23840 8870
rect 19550 8810 19770 8820
rect 19550 8610 19562 8810
rect 19762 8610 19770 8810
rect 19550 8600 19770 8610
rect 23520 8560 23530 8860
rect 23830 8560 23840 8860
rect 23520 8550 23840 8560
rect 25690 7720 25910 7730
rect 23060 7690 23200 7700
rect 21690 7660 21830 7670
rect 21690 7540 21700 7660
rect 21820 7540 21830 7660
rect 23060 7570 23070 7690
rect 23190 7570 23200 7690
rect 23060 7560 23200 7570
rect 21690 7530 21830 7540
rect 25690 7540 25710 7720
rect 25890 7540 25910 7720
rect 25690 7510 25910 7540
<< via2 >>
rect 25372 17112 25428 17168
rect 25932 16312 25988 16368
rect 25370 14440 25430 14500
rect 25930 14470 25990 14530
rect 19962 10290 20162 10490
rect 23485 10245 23775 10535
rect 19562 8610 19762 8810
rect 23535 8565 23825 8855
rect 21705 7545 21815 7655
rect 23075 7575 23185 7685
rect 25715 7545 25885 7715
<< metal3 >>
rect 25350 17172 25450 17190
rect 25350 17108 25368 17172
rect 25432 17108 25450 17172
rect 25350 17090 25450 17108
rect 25910 16372 26010 16390
rect 25910 16308 25928 16372
rect 25992 16308 26010 16372
rect 25910 16290 26010 16308
rect 681 16060 979 16065
rect 680 16059 16010 16060
rect 680 15761 681 16059
rect 979 15761 16010 16059
rect 680 15760 16010 15761
rect 681 15755 979 15760
rect 10297 15254 10595 15259
rect 10296 15253 15590 15254
rect 10296 14955 10297 15253
rect 10595 14955 15590 15253
rect 10296 14954 15590 14955
rect 10297 14949 10595 14954
rect 15480 14670 15590 14954
rect 15900 14650 16010 15760
rect 31283 15460 31461 15465
rect 16310 15459 31462 15460
rect 16310 15281 31283 15459
rect 31461 15281 31462 15459
rect 16310 15280 31462 15281
rect 16310 14510 16420 15280
rect 31283 15275 31461 15280
rect 16712 15048 16718 15112
rect 16782 15048 16788 15112
rect 16720 14580 16780 15048
rect 17512 15018 17518 15082
rect 17582 15018 17588 15082
rect 17128 14922 17192 14928
rect 17128 14852 17192 14858
rect 17130 14570 17190 14852
rect 17520 14590 17580 15018
rect 25925 14530 25995 14535
rect 25365 14500 25435 14505
rect 25365 14440 25370 14500
rect 25430 14440 25435 14500
rect 25925 14470 25930 14530
rect 25990 14470 25995 14530
rect 25925 14465 25995 14470
rect 25365 14435 25435 14440
rect 25370 12710 25430 14435
rect 25930 12730 25990 14465
rect 881 10540 1179 10545
rect 880 10539 23780 10540
rect 880 10241 881 10539
rect 1179 10535 23780 10539
rect 1179 10490 23485 10535
rect 1179 10290 19962 10490
rect 20162 10290 23485 10490
rect 1179 10245 23485 10290
rect 23775 10245 23780 10535
rect 1179 10241 23780 10245
rect 880 10240 23780 10241
rect 881 10235 1179 10240
rect 10501 8860 10799 8865
rect 10500 8859 23830 8860
rect 10500 8561 10501 8859
rect 10799 8855 23830 8859
rect 10799 8810 23535 8855
rect 10799 8610 19562 8810
rect 19762 8610 23535 8810
rect 10799 8565 23535 8610
rect 23825 8565 23830 8855
rect 10799 8561 23830 8565
rect 10500 8560 23830 8561
rect 10501 8555 10799 8560
rect 25358 8340 25478 8532
rect 21700 8220 25478 8340
rect 21700 7655 21820 8220
rect 25902 8080 26022 8532
rect 21700 7545 21705 7655
rect 21815 7545 21820 7655
rect 23070 7960 26022 8080
rect 23070 7685 23190 7960
rect 25711 7720 25889 7725
rect 23070 7575 23075 7685
rect 23185 7575 23190 7685
rect 23070 7570 23190 7575
rect 25710 7719 25890 7720
rect 21700 7540 21820 7545
rect 25710 7541 25711 7719
rect 25889 7541 25890 7719
rect 25710 7540 25890 7541
rect 25711 7535 25889 7540
<< via3 >>
rect 25368 17168 25432 17172
rect 25368 17112 25372 17168
rect 25372 17112 25428 17168
rect 25428 17112 25432 17168
rect 25368 17108 25432 17112
rect 25928 16368 25992 16372
rect 25928 16312 25932 16368
rect 25932 16312 25988 16368
rect 25988 16312 25992 16368
rect 25928 16308 25992 16312
rect 681 15761 979 16059
rect 10297 14955 10595 15253
rect 31283 15281 31461 15459
rect 16718 15048 16782 15112
rect 17518 15018 17582 15082
rect 17128 14858 17192 14922
rect 881 10241 1179 10539
rect 10501 8561 10799 8859
rect 25711 7715 25889 7719
rect 25711 7545 25715 7715
rect 25715 7545 25885 7715
rect 25885 7545 25889 7715
rect 25711 7541 25889 7545
<< metal4 >>
rect 798 44880 858 45152
rect 1534 44880 1594 45152
rect 2270 44880 2330 45152
rect 3006 44880 3066 45152
rect 3742 44880 3802 45152
rect 4478 44880 4538 45152
rect 5214 44880 5274 45152
rect 5950 44880 6010 45152
rect 6686 44880 6746 45152
rect 7422 44880 7482 45152
rect 8158 44880 8218 45152
rect 8894 44880 8954 45152
rect 9630 44880 9690 45152
rect 10366 44880 10426 45152
rect 11102 44880 11162 45152
rect 11838 44880 11898 45152
rect 12574 44880 12634 45152
rect 13310 44880 13370 45152
rect 14046 44880 14106 45152
rect 14782 44880 14842 45152
rect 15518 44880 15578 45152
rect 16254 44880 16314 45152
rect 16990 44880 17050 45152
rect 590 44570 17410 44880
rect 200 16060 500 44152
rect 200 16059 980 16060
rect 200 15761 681 16059
rect 979 15761 980 16059
rect 200 15760 980 15761
rect 200 10540 500 15760
rect 9800 15254 10100 44152
rect 17726 17250 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 16720 17190 17786 17250
rect 9800 15253 10596 15254
rect 9800 14955 10297 15253
rect 10595 14955 10596 15253
rect 16720 15113 16780 17190
rect 25367 17172 25433 17173
rect 25367 17108 25368 17172
rect 25432 17170 25433 17172
rect 27294 17170 27354 45152
rect 25432 17110 27354 17170
rect 25432 17108 25433 17110
rect 25367 17107 25433 17108
rect 25927 16372 25993 16373
rect 25927 16308 25928 16372
rect 25992 16370 25993 16372
rect 28030 16370 28090 45152
rect 25992 16310 28090 16370
rect 25992 16308 25993 16310
rect 25927 16307 25993 16308
rect 28766 15710 28826 45152
rect 17520 15650 28826 15710
rect 16717 15112 16783 15113
rect 16717 15048 16718 15112
rect 16782 15048 16783 15112
rect 17520 15083 17580 15650
rect 16717 15047 16783 15048
rect 17517 15082 17583 15083
rect 17517 15018 17518 15082
rect 17582 15018 17583 15082
rect 17517 15017 17583 15018
rect 9800 14954 10596 14955
rect 200 10539 1180 10540
rect 200 10241 881 10539
rect 1179 10241 1180 10539
rect 200 10240 1180 10241
rect 200 1000 500 10240
rect 9800 8860 10100 14954
rect 17127 14922 17193 14923
rect 17127 14858 17128 14922
rect 17192 14920 17193 14922
rect 29502 14920 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 17192 14860 29562 14920
rect 31282 15459 31462 15460
rect 31282 15281 31283 15459
rect 31461 15281 31462 15459
rect 17192 14858 17193 14860
rect 17127 14857 17193 14858
rect 9800 8859 10800 8860
rect 9800 8561 10501 8859
rect 10799 8561 10800 8859
rect 9800 8560 10800 8561
rect 9800 1000 10100 8560
rect 25710 7719 30600 7720
rect 25710 7541 25711 7719
rect 25889 7541 30600 7719
rect 25710 7540 30600 7541
rect 30420 3850 30600 7540
rect 26866 3670 30600 3850
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 3670
rect 31282 0 31462 15281
use charge_pump  charge_pump_0
timestamp 1717195371
transform 1 0 17712 0 1 5686
box 1850 -1570 12612 2030
use pfd  pfd_0
timestamp 1717194565
transform 0 1 25078 1 0 8412
box -38 -48 4400 1136
use vco  vco_0
timestamp 1717194565
transform 1 0 16000 0 1 12466
box -530 -1206 4600 2230
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
