magic
tech sky130A
magscale 1 2
timestamp 1717118324
<< viali >>
rect 2237 9605 2271 9639
rect 2881 9537 2915 9571
rect 857 9469 891 9503
rect 3433 9469 3467 9503
rect 3801 9469 3835 9503
rect 3893 9469 3927 9503
rect 4169 9469 4203 9503
rect 5917 9469 5951 9503
rect 6837 9469 6871 9503
rect 8401 9469 8435 9503
rect 1124 9401 1158 9435
rect 4414 9401 4448 9435
rect 7104 9401 7138 9435
rect 8646 9401 8680 9435
rect 2329 9333 2363 9367
rect 3249 9333 3283 9367
rect 3617 9333 3651 9367
rect 4077 9333 4111 9367
rect 5549 9333 5583 9367
rect 6561 9333 6595 9367
rect 8217 9333 8251 9367
rect 9781 9333 9815 9367
rect 1225 9129 1259 9163
rect 5641 9129 5675 9163
rect 3056 9061 3090 9095
rect 1041 8993 1075 9027
rect 1573 8993 1607 9027
rect 2789 8993 2823 9027
rect 4528 8993 4562 9027
rect 5917 8993 5951 9027
rect 6184 8993 6218 9027
rect 7389 8993 7423 9027
rect 7849 8993 7883 9027
rect 9873 8993 9907 9027
rect 1317 8925 1351 8959
rect 4261 8925 4295 8959
rect 9597 8925 9631 8959
rect 2697 8789 2731 8823
rect 4169 8789 4203 8823
rect 7297 8789 7331 8823
rect 7573 8789 7607 8823
rect 9689 8789 9723 8823
rect 1041 8585 1075 8619
rect 6561 8585 6595 8619
rect 6837 8585 6871 8619
rect 7941 8585 7975 8619
rect 8585 8517 8619 8551
rect 1685 8449 1719 8483
rect 5825 8449 5859 8483
rect 7757 8449 7791 8483
rect 857 8381 891 8415
rect 1409 8381 1443 8415
rect 5089 8381 5123 8415
rect 6745 8381 6779 8415
rect 7021 8381 7055 8415
rect 8125 8381 8159 8415
rect 9965 8381 9999 8415
rect 1930 8313 1964 8347
rect 3249 8313 3283 8347
rect 9698 8313 9732 8347
rect 1593 8245 1627 8279
rect 3065 8245 3099 8279
rect 4537 8245 4571 8279
rect 5733 8245 5767 8279
rect 6469 8245 6503 8279
rect 7205 8245 7239 8279
rect 4813 8041 4847 8075
rect 9781 8041 9815 8075
rect 1400 7973 1434 8007
rect 3678 7973 3712 8007
rect 1133 7905 1167 7939
rect 2697 7905 2731 7939
rect 5641 7905 5675 7939
rect 5825 7905 5859 7939
rect 6092 7905 6126 7939
rect 7389 7905 7423 7939
rect 7656 7905 7690 7939
rect 9597 7905 9631 7939
rect 3433 7837 3467 7871
rect 8861 7837 8895 7871
rect 2513 7701 2547 7735
rect 3341 7701 3375 7735
rect 4997 7701 5031 7735
rect 7205 7701 7239 7735
rect 8769 7701 8803 7735
rect 9505 7701 9539 7735
rect 8401 7497 8435 7531
rect 2789 7361 2823 7395
rect 3341 7361 3375 7395
rect 4169 7361 4203 7395
rect 6837 7361 6871 7395
rect 2053 7293 2087 7327
rect 2605 7293 2639 7327
rect 4905 7293 4939 7327
rect 5172 7293 5206 7327
rect 7104 7293 7138 7327
rect 9781 7293 9815 7327
rect 9514 7225 9548 7259
rect 1501 7157 1535 7191
rect 2421 7157 2455 7191
rect 3985 7157 4019 7191
rect 4813 7157 4847 7191
rect 6285 7157 6319 7191
rect 8217 7157 8251 7191
rect 3065 6885 3099 6919
rect 4436 6885 4470 6919
rect 9698 6885 9732 6919
rect 1225 6817 1259 6851
rect 1492 6817 1526 6851
rect 3525 6817 3559 6851
rect 4169 6817 4203 6851
rect 5825 6817 5859 6851
rect 6092 6817 6126 6851
rect 7941 6817 7975 6851
rect 8493 6817 8527 6851
rect 9965 6817 9999 6851
rect 3157 6749 3191 6783
rect 3249 6749 3283 6783
rect 2605 6681 2639 6715
rect 2697 6613 2731 6647
rect 3617 6613 3651 6647
rect 5549 6613 5583 6647
rect 7205 6613 7239 6647
rect 8585 6613 8619 6647
rect 3065 6409 3099 6443
rect 2329 6341 2363 6375
rect 4629 6341 4663 6375
rect 6745 6341 6779 6375
rect 2513 6273 2547 6307
rect 6101 6273 6135 6307
rect 7021 6273 7055 6307
rect 7297 6273 7331 6307
rect 7941 6273 7975 6307
rect 9781 6273 9815 6307
rect 949 6205 983 6239
rect 3249 6205 3283 6239
rect 3516 6205 3550 6239
rect 6285 6205 6319 6239
rect 7138 6205 7172 6239
rect 1216 6137 1250 6171
rect 9514 6137 9548 6171
rect 8401 6069 8435 6103
rect 1685 5865 1719 5899
rect 2145 5865 2179 5899
rect 4261 5865 4295 5899
rect 8309 5865 8343 5899
rect 9597 5865 9631 5899
rect 3148 5797 3182 5831
rect 5825 5797 5859 5831
rect 7573 5797 7607 5831
rect 2053 5729 2087 5763
rect 4537 5729 4571 5763
rect 7665 5729 7699 5763
rect 7941 5729 7975 5763
rect 8677 5729 8711 5763
rect 9873 5729 9907 5763
rect 2237 5661 2271 5695
rect 2881 5661 2915 5695
rect 4629 5661 4663 5695
rect 8769 5661 8803 5695
rect 8953 5661 8987 5695
rect 4905 5593 4939 5627
rect 7757 5525 7791 5559
rect 8033 5525 8067 5559
rect 9781 5525 9815 5559
rect 7205 5321 7239 5355
rect 7389 5321 7423 5355
rect 9965 5321 9999 5355
rect 1685 5253 1719 5287
rect 4353 5185 4387 5219
rect 4629 5185 4663 5219
rect 8401 5185 8435 5219
rect 8677 5185 8711 5219
rect 9321 5185 9355 5219
rect 2789 5117 2823 5151
rect 3433 5117 3467 5151
rect 4261 5117 4295 5151
rect 5733 5117 5767 5151
rect 5917 5117 5951 5151
rect 6009 5117 6043 5151
rect 6101 5117 6135 5151
rect 6285 5117 6319 5151
rect 6561 5117 6595 5151
rect 6709 5117 6743 5151
rect 7026 5117 7060 5151
rect 7297 5117 7331 5151
rect 7665 5117 7699 5151
rect 8769 5117 8803 5151
rect 1961 5049 1995 5083
rect 2145 5049 2179 5083
rect 3249 5049 3283 5083
rect 6837 5049 6871 5083
rect 6929 5049 6963 5083
rect 1501 4981 1535 5015
rect 3617 4981 3651 5015
rect 6469 4981 6503 5015
rect 7849 4981 7883 5015
rect 7757 4777 7791 4811
rect 1216 4709 1250 4743
rect 4537 4709 4571 4743
rect 8217 4709 8251 4743
rect 9781 4709 9815 4743
rect 2513 4641 2547 4675
rect 2697 4641 2731 4675
rect 4629 4641 4663 4675
rect 4813 4641 4847 4675
rect 5268 4641 5302 4675
rect 5365 4641 5399 4675
rect 5457 4641 5491 4675
rect 5641 4641 5675 4675
rect 6469 4641 6503 4675
rect 6653 4641 6687 4675
rect 6837 4641 6871 4675
rect 7021 4641 7055 4675
rect 7113 4641 7147 4675
rect 7261 4641 7295 4675
rect 7389 4641 7423 4675
rect 7481 4641 7515 4675
rect 7619 4641 7653 4675
rect 949 4573 983 4607
rect 6745 4573 6779 4607
rect 2329 4437 2363 4471
rect 2605 4437 2639 4471
rect 3249 4437 3283 4471
rect 4721 4437 4755 4471
rect 5641 4437 5675 4471
rect 6285 4437 6319 4471
rect 2697 4233 2731 4267
rect 3433 4233 3467 4267
rect 4997 4233 5031 4267
rect 6929 4233 6963 4267
rect 7481 4233 7515 4267
rect 8493 4233 8527 4267
rect 4261 4165 4295 4199
rect 6377 4165 6411 4199
rect 2973 4097 3007 4131
rect 5273 4097 5307 4131
rect 1317 4029 1351 4063
rect 2881 4029 2915 4063
rect 3065 4029 3099 4063
rect 3709 4029 3743 4063
rect 3893 4029 3927 4063
rect 4629 4029 4663 4063
rect 5089 4029 5123 4063
rect 5181 4029 5215 4063
rect 6561 4029 6595 4063
rect 7205 4029 7239 4063
rect 7297 4029 7331 4063
rect 7573 4029 7607 4063
rect 9873 4029 9907 4063
rect 1584 3961 1618 3995
rect 3417 3961 3451 3995
rect 3617 3961 3651 3995
rect 4537 3961 4571 3995
rect 6653 3961 6687 3995
rect 7021 3961 7055 3995
rect 9606 3961 9640 3995
rect 3249 3893 3283 3927
rect 4077 3893 4111 3927
rect 4445 3893 4479 3927
rect 4813 3893 4847 3927
rect 6745 3893 6779 3927
rect 3801 3689 3835 3723
rect 5273 3689 5307 3723
rect 7297 3689 7331 3723
rect 7665 3689 7699 3723
rect 9045 3689 9079 3723
rect 2421 3553 2455 3587
rect 2688 3553 2722 3587
rect 4160 3553 4194 3587
rect 7389 3553 7423 3587
rect 7757 3553 7791 3587
rect 7849 3553 7883 3587
rect 8033 3553 8067 3587
rect 8309 3553 8343 3587
rect 8401 3553 8435 3587
rect 8585 3553 8619 3587
rect 8677 3553 8711 3587
rect 8815 3553 8849 3587
rect 9137 3553 9171 3587
rect 9321 3553 9355 3587
rect 3893 3485 3927 3519
rect 7941 3417 7975 3451
rect 9505 3417 9539 3451
rect 8217 3349 8251 3383
rect 3249 3145 3283 3179
rect 3433 3145 3467 3179
rect 3985 3145 4019 3179
rect 4169 3145 4203 3179
rect 4537 3145 4571 3179
rect 8033 3145 8067 3179
rect 8493 3145 8527 3179
rect 7849 3077 7883 3111
rect 4629 2941 4663 2975
rect 7665 2941 7699 2975
rect 9873 2941 9907 2975
rect 3401 2873 3435 2907
rect 3617 2873 3651 2907
rect 4353 2873 4387 2907
rect 7481 2873 7515 2907
rect 8217 2873 8251 2907
rect 9606 2873 9640 2907
rect 4153 2805 4187 2839
rect 8017 2805 8051 2839
rect 6469 2601 6503 2635
rect 7481 2601 7515 2635
rect 8493 2601 8527 2635
rect 5441 2533 5475 2567
rect 5641 2533 5675 2567
rect 5825 2533 5859 2567
rect 6025 2533 6059 2567
rect 6653 2533 6687 2567
rect 7941 2533 7975 2567
rect 8125 2533 8159 2567
rect 8341 2533 8375 2567
rect 4721 2465 4755 2499
rect 4905 2465 4939 2499
rect 6561 2465 6595 2499
rect 6837 2465 6871 2499
rect 7205 2465 7239 2499
rect 7297 2465 7331 2499
rect 7481 2465 7515 2499
rect 7757 2465 7791 2499
rect 6285 2329 6319 2363
rect 4813 2261 4847 2295
rect 5273 2261 5307 2295
rect 5457 2261 5491 2295
rect 6009 2261 6043 2295
rect 6193 2261 6227 2295
rect 7113 2261 7147 2295
rect 7573 2261 7607 2295
rect 8309 2261 8343 2295
rect 4261 2057 4295 2091
rect 6377 2057 6411 2091
rect 6837 2057 6871 2091
rect 7113 2057 7147 2091
rect 7757 2057 7791 2091
rect 8401 2057 8435 2091
rect 4997 1921 5031 1955
rect 4905 1853 4939 1887
rect 5264 1853 5298 1887
rect 6469 1853 6503 1887
rect 6653 1853 6687 1887
rect 9781 1853 9815 1887
rect 4077 1785 4111 1819
rect 4293 1785 4327 1819
rect 4537 1785 4571 1819
rect 4721 1785 4755 1819
rect 7097 1785 7131 1819
rect 7297 1785 7331 1819
rect 7573 1785 7607 1819
rect 7789 1785 7823 1819
rect 9514 1785 9548 1819
rect 4445 1717 4479 1751
rect 6929 1717 6963 1751
rect 7941 1717 7975 1751
rect 6469 1513 6503 1547
rect 6837 1513 6871 1547
rect 4517 1445 4551 1479
rect 7950 1445 7984 1479
rect 4261 1377 4295 1411
rect 6009 1377 6043 1411
rect 6193 1377 6227 1411
rect 6285 1377 6319 1411
rect 6377 1377 6411 1411
rect 5825 1309 5859 1343
rect 8217 1309 8251 1343
rect 5641 1241 5675 1275
rect 2789 901 2823 935
rect 8585 901 8619 935
rect 2973 765 3007 799
rect 8401 765 8435 799
<< metal1 >>
rect 552 9818 10304 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 10304 9818
rect 552 9744 10304 9766
rect 4522 9704 4528 9716
rect 3896 9676 4528 9704
rect 2225 9639 2283 9645
rect 2225 9605 2237 9639
rect 2271 9636 2283 9639
rect 2271 9608 2774 9636
rect 2271 9605 2283 9608
rect 2225 9599 2283 9605
rect 2746 9568 2774 9608
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 2746 9540 2881 9568
rect 2869 9537 2881 9540
rect 2915 9537 2927 9571
rect 2869 9531 2927 9537
rect 845 9503 903 9509
rect 845 9469 857 9503
rect 891 9500 903 9503
rect 891 9472 1256 9500
rect 891 9469 903 9472
rect 845 9463 903 9469
rect 1228 9444 1256 9472
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 3421 9503 3479 9509
rect 3421 9500 3433 9503
rect 3016 9472 3433 9500
rect 3016 9460 3022 9472
rect 3421 9469 3433 9472
rect 3467 9469 3479 9503
rect 3421 9463 3479 9469
rect 3510 9460 3516 9512
rect 3568 9500 3574 9512
rect 3896 9509 3924 9676
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 3789 9503 3847 9509
rect 3789 9500 3801 9503
rect 3568 9472 3801 9500
rect 3568 9460 3574 9472
rect 3789 9469 3801 9472
rect 3835 9469 3847 9503
rect 3789 9463 3847 9469
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 4154 9460 4160 9512
rect 4212 9460 4218 9512
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 5905 9503 5963 9509
rect 5905 9500 5917 9503
rect 5684 9472 5917 9500
rect 5684 9460 5690 9472
rect 5905 9469 5917 9472
rect 5951 9469 5963 9503
rect 5905 9463 5963 9469
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 6880 9472 8401 9500
rect 6880 9460 6886 9472
rect 8389 9469 8401 9472
rect 8435 9500 8447 9503
rect 9950 9500 9956 9512
rect 8435 9472 9956 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 9950 9460 9956 9472
rect 10008 9460 10014 9512
rect 1118 9441 1124 9444
rect 1112 9395 1124 9441
rect 1118 9392 1124 9395
rect 1176 9392 1182 9444
rect 1210 9392 1216 9444
rect 1268 9392 1274 9444
rect 4402 9435 4460 9441
rect 4402 9432 4414 9435
rect 4080 9404 4414 9432
rect 2314 9324 2320 9376
rect 2372 9324 2378 9376
rect 3234 9324 3240 9376
rect 3292 9324 3298 9376
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 4080 9373 4108 9404
rect 4402 9401 4414 9404
rect 4448 9401 4460 9435
rect 4402 9395 4460 9401
rect 7092 9435 7150 9441
rect 7092 9401 7104 9435
rect 7138 9432 7150 9435
rect 7742 9432 7748 9444
rect 7138 9404 7748 9432
rect 7138 9401 7150 9404
rect 7092 9395 7150 9401
rect 7742 9392 7748 9404
rect 7800 9392 7806 9444
rect 7852 9404 8340 9432
rect 3605 9367 3663 9373
rect 3605 9364 3617 9367
rect 3568 9336 3617 9364
rect 3568 9324 3574 9336
rect 3605 9333 3617 9336
rect 3651 9333 3663 9367
rect 3605 9327 3663 9333
rect 4065 9367 4123 9373
rect 4065 9333 4077 9367
rect 4111 9333 4123 9367
rect 4065 9327 4123 9333
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 5810 9364 5816 9376
rect 5583 9336 5816 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 6546 9324 6552 9376
rect 6604 9324 6610 9376
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 7852 9364 7880 9404
rect 7432 9336 7880 9364
rect 7432 9324 7438 9336
rect 8110 9324 8116 9376
rect 8168 9364 8174 9376
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 8168 9336 8217 9364
rect 8168 9324 8174 9336
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 8312 9364 8340 9404
rect 8478 9392 8484 9444
rect 8536 9432 8542 9444
rect 8634 9435 8692 9441
rect 8634 9432 8646 9435
rect 8536 9404 8646 9432
rect 8536 9392 8542 9404
rect 8634 9401 8646 9404
rect 8680 9401 8692 9435
rect 8634 9395 8692 9401
rect 9769 9367 9827 9373
rect 9769 9364 9781 9367
rect 8312 9336 9781 9364
rect 8205 9327 8263 9333
rect 9769 9333 9781 9336
rect 9815 9333 9827 9367
rect 9769 9327 9827 9333
rect 552 9274 10304 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 10304 9274
rect 552 9200 10304 9222
rect 1213 9163 1271 9169
rect 1213 9129 1225 9163
rect 1259 9129 1271 9163
rect 1213 9123 1271 9129
rect 1026 8984 1032 9036
rect 1084 8984 1090 9036
rect 1228 9024 1256 9123
rect 5626 9120 5632 9172
rect 5684 9120 5690 9172
rect 3044 9095 3102 9101
rect 3044 9061 3056 9095
rect 3090 9092 3102 9095
rect 3234 9092 3240 9104
rect 3090 9064 3240 9092
rect 3090 9061 3102 9064
rect 3044 9055 3102 9061
rect 3234 9052 3240 9064
rect 3292 9052 3298 9104
rect 6822 9092 6828 9104
rect 5920 9064 6828 9092
rect 1561 9027 1619 9033
rect 1561 9024 1573 9027
rect 1228 8996 1573 9024
rect 1561 8993 1573 8996
rect 1607 8993 1619 9027
rect 2777 9027 2835 9033
rect 2777 9024 2789 9027
rect 1561 8987 1619 8993
rect 2332 8996 2789 9024
rect 1210 8916 1216 8968
rect 1268 8956 1274 8968
rect 1305 8959 1363 8965
rect 1305 8956 1317 8959
rect 1268 8928 1317 8956
rect 1268 8916 1274 8928
rect 1305 8925 1317 8928
rect 1351 8925 1363 8959
rect 1305 8919 1363 8925
rect 1320 8820 1348 8919
rect 2332 8820 2360 8996
rect 2777 8993 2789 8996
rect 2823 8993 2835 9027
rect 2777 8987 2835 8993
rect 4516 9027 4574 9033
rect 4516 8993 4528 9027
rect 4562 9024 4574 9027
rect 5718 9024 5724 9036
rect 4562 8996 5724 9024
rect 4562 8993 4574 8996
rect 4516 8987 4574 8993
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 5920 9033 5948 9064
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 6172 9027 6230 9033
rect 6172 8993 6184 9027
rect 6218 9024 6230 9027
rect 6730 9024 6736 9036
rect 6218 8996 6736 9024
rect 6218 8993 6230 8996
rect 6172 8987 6230 8993
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 7006 8984 7012 9036
rect 7064 9024 7070 9036
rect 7377 9027 7435 9033
rect 7377 9024 7389 9027
rect 7064 8996 7389 9024
rect 7064 8984 7070 8996
rect 7377 8993 7389 8996
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 7834 8984 7840 9036
rect 7892 8984 7898 9036
rect 8662 8984 8668 9036
rect 8720 9024 8726 9036
rect 9861 9027 9919 9033
rect 9861 9024 9873 9027
rect 8720 8996 9873 9024
rect 8720 8984 8726 8996
rect 9861 8993 9873 8996
rect 9907 8993 9919 9027
rect 9861 8987 9919 8993
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 4249 8959 4307 8965
rect 4249 8956 4261 8959
rect 4212 8928 4261 8956
rect 4212 8916 4218 8928
rect 4249 8925 4261 8928
rect 4295 8925 4307 8959
rect 4249 8919 4307 8925
rect 9585 8959 9643 8965
rect 9585 8925 9597 8959
rect 9631 8956 9643 8959
rect 9950 8956 9956 8968
rect 9631 8928 9956 8956
rect 9631 8925 9643 8928
rect 9585 8919 9643 8925
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 1320 8792 2360 8820
rect 2682 8780 2688 8832
rect 2740 8780 2746 8832
rect 4157 8823 4215 8829
rect 4157 8789 4169 8823
rect 4203 8820 4215 8823
rect 4246 8820 4252 8832
rect 4203 8792 4252 8820
rect 4203 8789 4215 8792
rect 4157 8783 4215 8789
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 7282 8780 7288 8832
rect 7340 8780 7346 8832
rect 7561 8823 7619 8829
rect 7561 8789 7573 8823
rect 7607 8820 7619 8823
rect 7650 8820 7656 8832
rect 7607 8792 7656 8820
rect 7607 8789 7619 8792
rect 7561 8783 7619 8789
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 9398 8780 9404 8832
rect 9456 8820 9462 8832
rect 9677 8823 9735 8829
rect 9677 8820 9689 8823
rect 9456 8792 9689 8820
rect 9456 8780 9462 8792
rect 9677 8789 9689 8792
rect 9723 8789 9735 8823
rect 9677 8783 9735 8789
rect 552 8730 10304 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 10304 8730
rect 552 8656 10304 8678
rect 1029 8619 1087 8625
rect 1029 8585 1041 8619
rect 1075 8616 1087 8619
rect 1118 8616 1124 8628
rect 1075 8588 1124 8616
rect 1075 8585 1087 8588
rect 1029 8579 1087 8585
rect 1118 8576 1124 8588
rect 1176 8576 1182 8628
rect 5718 8576 5724 8628
rect 5776 8616 5782 8628
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 5776 8588 6561 8616
rect 5776 8576 5782 8588
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 6549 8579 6607 8585
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 6788 8588 6837 8616
rect 6788 8576 6794 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 6825 8579 6883 8585
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 7929 8619 7987 8625
rect 7929 8616 7941 8619
rect 7800 8588 7941 8616
rect 7800 8576 7806 8588
rect 7929 8585 7941 8588
rect 7975 8585 7987 8619
rect 7929 8579 7987 8585
rect 5626 8508 5632 8560
rect 5684 8548 5690 8560
rect 8573 8551 8631 8557
rect 8573 8548 8585 8551
rect 5684 8520 8585 8548
rect 5684 8508 5690 8520
rect 8573 8517 8585 8520
rect 8619 8517 8631 8551
rect 8573 8511 8631 8517
rect 1210 8440 1216 8492
rect 1268 8480 1274 8492
rect 1673 8483 1731 8489
rect 1673 8480 1685 8483
rect 1268 8452 1685 8480
rect 1268 8440 1274 8452
rect 1673 8449 1685 8452
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 6178 8440 6184 8492
rect 6236 8480 6242 8492
rect 6236 8452 7052 8480
rect 6236 8440 6242 8452
rect 382 8372 388 8424
rect 440 8412 446 8424
rect 845 8415 903 8421
rect 845 8412 857 8415
rect 440 8384 857 8412
rect 440 8372 446 8384
rect 845 8381 857 8384
rect 891 8381 903 8415
rect 845 8375 903 8381
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1443 8384 2084 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2056 8356 2084 8384
rect 5074 8372 5080 8424
rect 5132 8372 5138 8424
rect 5350 8372 5356 8424
rect 5408 8412 5414 8424
rect 7024 8421 7052 8452
rect 7282 8440 7288 8492
rect 7340 8480 7346 8492
rect 7745 8483 7803 8489
rect 7745 8480 7757 8483
rect 7340 8452 7757 8480
rect 7340 8440 7346 8452
rect 7745 8449 7757 8452
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 6733 8415 6791 8421
rect 6733 8412 6745 8415
rect 5408 8384 6745 8412
rect 5408 8372 5414 8384
rect 6733 8381 6745 8384
rect 6779 8381 6791 8415
rect 6733 8375 6791 8381
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8381 7067 8415
rect 7009 8375 7067 8381
rect 7926 8372 7932 8424
rect 7984 8412 7990 8424
rect 8113 8415 8171 8421
rect 8113 8412 8125 8415
rect 7984 8384 8125 8412
rect 7984 8372 7990 8384
rect 8113 8381 8125 8384
rect 8159 8381 8171 8415
rect 8113 8375 8171 8381
rect 9950 8372 9956 8424
rect 10008 8372 10014 8424
rect 1918 8347 1976 8353
rect 1918 8344 1930 8347
rect 1596 8316 1930 8344
rect 1596 8285 1624 8316
rect 1918 8313 1930 8316
rect 1964 8313 1976 8347
rect 1918 8307 1976 8313
rect 2038 8304 2044 8356
rect 2096 8304 2102 8356
rect 3237 8347 3295 8353
rect 3237 8313 3249 8347
rect 3283 8344 3295 8347
rect 5534 8344 5540 8356
rect 3283 8316 5540 8344
rect 3283 8313 3295 8316
rect 3237 8307 3295 8313
rect 5534 8304 5540 8316
rect 5592 8344 5598 8356
rect 7834 8344 7840 8356
rect 5592 8316 7840 8344
rect 5592 8304 5598 8316
rect 7834 8304 7840 8316
rect 7892 8304 7898 8356
rect 9674 8304 9680 8356
rect 9732 8353 9738 8356
rect 9732 8307 9744 8353
rect 9732 8304 9738 8307
rect 1581 8279 1639 8285
rect 1581 8245 1593 8279
rect 1627 8245 1639 8279
rect 1581 8239 1639 8245
rect 3050 8236 3056 8288
rect 3108 8236 3114 8288
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4525 8279 4583 8285
rect 4525 8276 4537 8279
rect 4212 8248 4537 8276
rect 4212 8236 4218 8248
rect 4525 8245 4537 8248
rect 4571 8245 4583 8279
rect 4525 8239 4583 8245
rect 5718 8236 5724 8288
rect 5776 8236 5782 8288
rect 6454 8236 6460 8288
rect 6512 8236 6518 8288
rect 7098 8236 7104 8288
rect 7156 8276 7162 8288
rect 7193 8279 7251 8285
rect 7193 8276 7205 8279
rect 7156 8248 7205 8276
rect 7156 8236 7162 8248
rect 7193 8245 7205 8248
rect 7239 8245 7251 8279
rect 7193 8239 7251 8245
rect 552 8186 10304 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 10304 8186
rect 552 8112 10304 8134
rect 4801 8075 4859 8081
rect 4801 8041 4813 8075
rect 4847 8072 4859 8075
rect 5074 8072 5080 8084
rect 4847 8044 5080 8072
rect 4847 8041 4859 8044
rect 4801 8035 4859 8041
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 9769 8075 9827 8081
rect 9769 8072 9781 8075
rect 9732 8044 9781 8072
rect 9732 8032 9738 8044
rect 9769 8041 9781 8044
rect 9815 8041 9827 8075
rect 9769 8035 9827 8041
rect 1388 8007 1446 8013
rect 1388 7973 1400 8007
rect 1434 8004 1446 8007
rect 2314 8004 2320 8016
rect 1434 7976 2320 8004
rect 1434 7973 1446 7976
rect 1388 7967 1446 7973
rect 2314 7964 2320 7976
rect 2372 7964 2378 8016
rect 3510 7964 3516 8016
rect 3568 8004 3574 8016
rect 3666 8007 3724 8013
rect 3666 8004 3678 8007
rect 3568 7976 3678 8004
rect 3568 7964 3574 7976
rect 3666 7973 3678 7976
rect 3712 7973 3724 8007
rect 3666 7967 3724 7973
rect 5828 7976 6868 8004
rect 1121 7939 1179 7945
rect 1121 7905 1133 7939
rect 1167 7936 1179 7939
rect 1210 7936 1216 7948
rect 1167 7908 1216 7936
rect 1167 7905 1179 7908
rect 1121 7899 1179 7905
rect 1210 7896 1216 7908
rect 1268 7896 1274 7948
rect 2682 7896 2688 7948
rect 2740 7896 2746 7948
rect 4154 7936 4160 7948
rect 3436 7908 4160 7936
rect 3436 7877 3464 7908
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 5626 7896 5632 7948
rect 5684 7896 5690 7948
rect 5828 7945 5856 7976
rect 6840 7948 6868 7976
rect 5813 7939 5871 7945
rect 5813 7905 5825 7939
rect 5859 7905 5871 7939
rect 5813 7899 5871 7905
rect 6080 7939 6138 7945
rect 6080 7905 6092 7939
rect 6126 7936 6138 7939
rect 6546 7936 6552 7948
rect 6126 7908 6552 7936
rect 6126 7905 6138 7908
rect 6080 7899 6138 7905
rect 6546 7896 6552 7908
rect 6604 7896 6610 7948
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 7650 7945 7656 7948
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 6880 7908 7389 7936
rect 6880 7896 6886 7908
rect 7377 7905 7389 7908
rect 7423 7905 7435 7939
rect 7644 7936 7656 7945
rect 7611 7908 7656 7936
rect 7377 7899 7435 7905
rect 7644 7899 7656 7908
rect 7650 7896 7656 7899
rect 7708 7896 7714 7948
rect 9490 7896 9496 7948
rect 9548 7936 9554 7948
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 9548 7908 9597 7936
rect 9548 7896 9554 7908
rect 9585 7905 9597 7908
rect 9631 7905 9643 7939
rect 9585 7899 9643 7905
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 8849 7871 8907 7877
rect 8849 7868 8861 7871
rect 8444 7840 8861 7868
rect 8444 7828 8450 7840
rect 8849 7837 8861 7840
rect 8895 7837 8907 7871
rect 8849 7831 8907 7837
rect 2501 7735 2559 7741
rect 2501 7701 2513 7735
rect 2547 7732 2559 7735
rect 2774 7732 2780 7744
rect 2547 7704 2780 7732
rect 2547 7701 2559 7704
rect 2501 7695 2559 7701
rect 2774 7692 2780 7704
rect 2832 7692 2838 7744
rect 3326 7692 3332 7744
rect 3384 7692 3390 7744
rect 4982 7692 4988 7744
rect 5040 7692 5046 7744
rect 7193 7735 7251 7741
rect 7193 7701 7205 7735
rect 7239 7732 7251 7735
rect 7282 7732 7288 7744
rect 7239 7704 7288 7732
rect 7239 7701 7251 7704
rect 7193 7695 7251 7701
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 8757 7735 8815 7741
rect 8757 7732 8769 7735
rect 8076 7704 8769 7732
rect 8076 7692 8082 7704
rect 8757 7701 8769 7704
rect 8803 7701 8815 7735
rect 8757 7695 8815 7701
rect 9490 7692 9496 7744
rect 9548 7692 9554 7744
rect 552 7642 10304 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 10304 7642
rect 552 7568 10304 7590
rect 8386 7488 8392 7540
rect 8444 7488 8450 7540
rect 4246 7460 4252 7472
rect 4172 7432 4252 7460
rect 2774 7352 2780 7404
rect 2832 7352 2838 7404
rect 3050 7352 3056 7404
rect 3108 7392 3114 7404
rect 4172 7401 4200 7432
rect 4246 7420 4252 7432
rect 4304 7420 4310 7472
rect 3329 7395 3387 7401
rect 3329 7392 3341 7395
rect 3108 7364 3341 7392
rect 3108 7352 3114 7364
rect 3329 7361 3341 7364
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 6822 7352 6828 7404
rect 6880 7352 6886 7404
rect 2038 7284 2044 7336
rect 2096 7284 2102 7336
rect 2498 7284 2504 7336
rect 2556 7324 2562 7336
rect 2593 7327 2651 7333
rect 2593 7324 2605 7327
rect 2556 7296 2605 7324
rect 2556 7284 2562 7296
rect 2593 7293 2605 7296
rect 2639 7293 2651 7327
rect 2593 7287 2651 7293
rect 4246 7284 4252 7336
rect 4304 7324 4310 7336
rect 4893 7327 4951 7333
rect 4893 7324 4905 7327
rect 4304 7296 4905 7324
rect 4304 7284 4310 7296
rect 4893 7293 4905 7296
rect 4939 7293 4951 7327
rect 4893 7287 4951 7293
rect 5160 7327 5218 7333
rect 5160 7293 5172 7327
rect 5206 7324 5218 7327
rect 5718 7324 5724 7336
rect 5206 7296 5724 7324
rect 5206 7293 5218 7296
rect 5160 7287 5218 7293
rect 5718 7284 5724 7296
rect 5776 7284 5782 7336
rect 7098 7333 7104 7336
rect 7092 7324 7104 7333
rect 7059 7296 7104 7324
rect 7092 7287 7104 7296
rect 7098 7284 7104 7287
rect 7156 7284 7162 7336
rect 9766 7284 9772 7336
rect 9824 7284 9830 7336
rect 9398 7216 9404 7268
rect 9456 7256 9462 7268
rect 9502 7259 9560 7265
rect 9502 7256 9514 7259
rect 9456 7228 9514 7256
rect 9456 7216 9462 7228
rect 9502 7225 9514 7228
rect 9548 7225 9560 7259
rect 9502 7219 9560 7225
rect 1302 7148 1308 7200
rect 1360 7188 1366 7200
rect 1489 7191 1547 7197
rect 1489 7188 1501 7191
rect 1360 7160 1501 7188
rect 1360 7148 1366 7160
rect 1489 7157 1501 7160
rect 1535 7157 1547 7191
rect 1489 7151 1547 7157
rect 2406 7148 2412 7200
rect 2464 7148 2470 7200
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 3973 7191 4031 7197
rect 3973 7188 3985 7191
rect 3568 7160 3985 7188
rect 3568 7148 3574 7160
rect 3973 7157 3985 7160
rect 4019 7157 4031 7191
rect 3973 7151 4031 7157
rect 4798 7148 4804 7200
rect 4856 7148 4862 7200
rect 6273 7191 6331 7197
rect 6273 7157 6285 7191
rect 6319 7188 6331 7191
rect 7006 7188 7012 7200
rect 6319 7160 7012 7188
rect 6319 7157 6331 7160
rect 6273 7151 6331 7157
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 8202 7148 8208 7200
rect 8260 7148 8266 7200
rect 552 7098 10304 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 10304 7098
rect 552 7024 10304 7046
rect 3053 6919 3111 6925
rect 3053 6916 3065 6919
rect 1228 6888 3065 6916
rect 1228 6860 1256 6888
rect 3053 6885 3065 6888
rect 3099 6916 3111 6919
rect 4424 6919 4482 6925
rect 3099 6888 4108 6916
rect 3099 6885 3111 6888
rect 3053 6879 3111 6885
rect 1210 6848 1216 6860
rect 1191 6820 1216 6848
rect 1210 6808 1216 6820
rect 1268 6808 1274 6860
rect 1480 6851 1538 6857
rect 1480 6817 1492 6851
rect 1526 6848 1538 6851
rect 1526 6820 3372 6848
rect 1526 6817 1538 6820
rect 1480 6811 1538 6817
rect 2498 6740 2504 6792
rect 2556 6780 2562 6792
rect 3145 6783 3203 6789
rect 3145 6780 3157 6783
rect 2556 6752 3157 6780
rect 2556 6740 2562 6752
rect 3145 6749 3157 6752
rect 3191 6749 3203 6783
rect 3145 6743 3203 6749
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6749 3295 6783
rect 3344 6780 3372 6820
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 3513 6851 3571 6857
rect 3513 6848 3525 6851
rect 3476 6820 3525 6848
rect 3476 6808 3482 6820
rect 3513 6817 3525 6820
rect 3559 6817 3571 6851
rect 4080 6848 4108 6888
rect 4424 6885 4436 6919
rect 4470 6916 4482 6919
rect 4798 6916 4804 6928
rect 4470 6888 4804 6916
rect 4470 6885 4482 6888
rect 4424 6879 4482 6885
rect 4798 6876 4804 6888
rect 4856 6876 4862 6928
rect 6822 6916 6828 6928
rect 5828 6888 6828 6916
rect 4154 6848 4160 6860
rect 4080 6820 4160 6848
rect 3513 6811 3571 6817
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 4982 6848 4988 6860
rect 4264 6820 4988 6848
rect 4264 6780 4292 6820
rect 4982 6808 4988 6820
rect 5040 6808 5046 6860
rect 5828 6857 5856 6888
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 9490 6876 9496 6928
rect 9548 6916 9554 6928
rect 9686 6919 9744 6925
rect 9686 6916 9698 6919
rect 9548 6888 9698 6916
rect 9548 6876 9554 6888
rect 9686 6885 9698 6888
rect 9732 6885 9744 6919
rect 9686 6879 9744 6885
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6817 5871 6851
rect 5813 6811 5871 6817
rect 6080 6851 6138 6857
rect 6080 6817 6092 6851
rect 6126 6848 6138 6851
rect 6454 6848 6460 6860
rect 6126 6820 6460 6848
rect 6126 6817 6138 6820
rect 6080 6811 6138 6817
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 7929 6851 7987 6857
rect 7929 6817 7941 6851
rect 7975 6848 7987 6851
rect 8018 6848 8024 6860
rect 7975 6820 8024 6848
rect 7975 6817 7987 6820
rect 7929 6811 7987 6817
rect 8018 6808 8024 6820
rect 8076 6808 8082 6860
rect 8478 6808 8484 6860
rect 8536 6808 8542 6860
rect 9950 6808 9956 6860
rect 10008 6808 10014 6860
rect 3344 6752 4292 6780
rect 3237 6743 3295 6749
rect 2593 6715 2651 6721
rect 2593 6681 2605 6715
rect 2639 6712 2651 6715
rect 3252 6712 3280 6743
rect 2639 6684 3280 6712
rect 2639 6681 2651 6684
rect 2593 6675 2651 6681
rect 2685 6647 2743 6653
rect 2685 6613 2697 6647
rect 2731 6644 2743 6647
rect 2958 6644 2964 6656
rect 2731 6616 2964 6644
rect 2731 6613 2743 6616
rect 2685 6607 2743 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 3050 6604 3056 6656
rect 3108 6644 3114 6656
rect 3605 6647 3663 6653
rect 3605 6644 3617 6647
rect 3108 6616 3617 6644
rect 3108 6604 3114 6616
rect 3605 6613 3617 6616
rect 3651 6613 3663 6647
rect 3605 6607 3663 6613
rect 5537 6647 5595 6653
rect 5537 6613 5549 6647
rect 5583 6644 5595 6647
rect 6086 6644 6092 6656
rect 5583 6616 6092 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 6086 6604 6092 6616
rect 6144 6644 6150 6656
rect 7098 6644 7104 6656
rect 6144 6616 7104 6644
rect 6144 6604 6150 6616
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7193 6647 7251 6653
rect 7193 6613 7205 6647
rect 7239 6644 7251 6647
rect 7926 6644 7932 6656
rect 7239 6616 7932 6644
rect 7239 6613 7251 6616
rect 7193 6607 7251 6613
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 8662 6644 8668 6656
rect 8619 6616 8668 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 8662 6604 8668 6616
rect 8720 6604 8726 6656
rect 552 6554 10304 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 10304 6554
rect 552 6480 10304 6502
rect 3053 6443 3111 6449
rect 3053 6409 3065 6443
rect 3099 6440 3111 6443
rect 3418 6440 3424 6452
rect 3099 6412 3424 6440
rect 3099 6409 3111 6412
rect 3053 6403 3111 6409
rect 3418 6400 3424 6412
rect 3476 6400 3482 6452
rect 7926 6440 7932 6452
rect 6748 6412 7932 6440
rect 6748 6381 6776 6412
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 2317 6375 2375 6381
rect 2317 6341 2329 6375
rect 2363 6341 2375 6375
rect 2317 6335 2375 6341
rect 4617 6375 4675 6381
rect 4617 6341 4629 6375
rect 4663 6341 4675 6375
rect 4617 6335 4675 6341
rect 6733 6375 6791 6381
rect 6733 6341 6745 6375
rect 6779 6341 6791 6375
rect 6733 6335 6791 6341
rect 2332 6304 2360 6335
rect 2498 6304 2504 6316
rect 2332 6276 2504 6304
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 4632 6304 4660 6335
rect 4706 6304 4712 6316
rect 4632 6276 4712 6304
rect 4706 6264 4712 6276
rect 4764 6304 4770 6316
rect 6089 6307 6147 6313
rect 6089 6304 6101 6307
rect 4764 6276 6101 6304
rect 4764 6264 4770 6276
rect 6089 6273 6101 6276
rect 6135 6273 6147 6307
rect 6089 6267 6147 6273
rect 7006 6264 7012 6316
rect 7064 6264 7070 6316
rect 7282 6264 7288 6316
rect 7340 6264 7346 6316
rect 7650 6264 7656 6316
rect 7708 6304 7714 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7708 6276 7941 6304
rect 7708 6264 7714 6276
rect 7929 6273 7941 6276
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 9766 6264 9772 6316
rect 9824 6264 9830 6316
rect 934 6196 940 6248
rect 992 6196 998 6248
rect 3234 6196 3240 6248
rect 3292 6196 3298 6248
rect 3510 6245 3516 6248
rect 3504 6236 3516 6245
rect 3471 6208 3516 6236
rect 3504 6199 3516 6208
rect 3510 6196 3516 6199
rect 3568 6196 3574 6248
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 6273 6239 6331 6245
rect 6273 6236 6285 6239
rect 4304 6208 6285 6236
rect 4304 6196 4310 6208
rect 6273 6205 6285 6208
rect 6319 6205 6331 6239
rect 6273 6199 6331 6205
rect 7098 6196 7104 6248
rect 7156 6245 7162 6248
rect 7156 6239 7184 6245
rect 7172 6205 7184 6239
rect 7156 6199 7184 6205
rect 7156 6196 7162 6199
rect 1204 6171 1262 6177
rect 1204 6137 1216 6171
rect 1250 6168 1262 6171
rect 1302 6168 1308 6180
rect 1250 6140 1308 6168
rect 1250 6137 1262 6140
rect 1204 6131 1262 6137
rect 1302 6128 1308 6140
rect 1360 6128 1366 6180
rect 9490 6128 9496 6180
rect 9548 6177 9554 6180
rect 9548 6131 9560 6177
rect 9548 6128 9554 6131
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 8389 6103 8447 6109
rect 8389 6100 8401 6103
rect 7156 6072 8401 6100
rect 7156 6060 7162 6072
rect 8389 6069 8401 6072
rect 8435 6069 8447 6103
rect 8389 6063 8447 6069
rect 552 6010 10304 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 10304 6010
rect 552 5936 10304 5958
rect 1673 5899 1731 5905
rect 1673 5865 1685 5899
rect 1719 5896 1731 5899
rect 2038 5896 2044 5908
rect 1719 5868 2044 5896
rect 1719 5865 1731 5868
rect 1673 5859 1731 5865
rect 2038 5856 2044 5868
rect 2096 5856 2102 5908
rect 2133 5899 2191 5905
rect 2133 5865 2145 5899
rect 2179 5896 2191 5899
rect 2406 5896 2412 5908
rect 2179 5868 2412 5896
rect 2179 5865 2191 5868
rect 2133 5859 2191 5865
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 3050 5896 3056 5908
rect 2746 5868 3056 5896
rect 2041 5763 2099 5769
rect 2041 5729 2053 5763
rect 2087 5760 2099 5763
rect 2746 5760 2774 5868
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 4246 5856 4252 5908
rect 4304 5856 4310 5908
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 8297 5899 8355 5905
rect 8297 5896 8309 5899
rect 7892 5868 8309 5896
rect 7892 5856 7898 5868
rect 8297 5865 8309 5868
rect 8343 5865 8355 5899
rect 8297 5859 8355 5865
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 9585 5899 9643 5905
rect 9585 5896 9597 5899
rect 9548 5868 9597 5896
rect 9548 5856 9554 5868
rect 9585 5865 9597 5868
rect 9631 5865 9643 5899
rect 9585 5859 9643 5865
rect 3136 5831 3194 5837
rect 3136 5797 3148 5831
rect 3182 5828 3194 5831
rect 3326 5828 3332 5840
rect 3182 5800 3332 5828
rect 3182 5797 3194 5800
rect 3136 5791 3194 5797
rect 3326 5788 3332 5800
rect 3384 5788 3390 5840
rect 5534 5788 5540 5840
rect 5592 5828 5598 5840
rect 5813 5831 5871 5837
rect 5813 5828 5825 5831
rect 5592 5800 5825 5828
rect 5592 5788 5598 5800
rect 5813 5797 5825 5800
rect 5859 5828 5871 5831
rect 7466 5828 7472 5840
rect 5859 5800 7472 5828
rect 5859 5797 5871 5800
rect 5813 5791 5871 5797
rect 7466 5788 7472 5800
rect 7524 5788 7530 5840
rect 7561 5831 7619 5837
rect 7561 5797 7573 5831
rect 7607 5828 7619 5831
rect 10318 5828 10324 5840
rect 7607 5800 10324 5828
rect 7607 5797 7619 5800
rect 7561 5791 7619 5797
rect 10318 5788 10324 5800
rect 10376 5788 10382 5840
rect 2087 5732 2774 5760
rect 2087 5729 2099 5732
rect 2041 5723 2099 5729
rect 4522 5720 4528 5772
rect 4580 5720 4586 5772
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 7340 5732 7665 5760
rect 7340 5720 7346 5732
rect 7653 5729 7665 5732
rect 7699 5729 7711 5763
rect 7653 5723 7711 5729
rect 7926 5720 7932 5772
rect 7984 5720 7990 5772
rect 8662 5720 8668 5772
rect 8720 5720 8726 5772
rect 9858 5720 9864 5772
rect 9916 5720 9922 5772
rect 2222 5652 2228 5704
rect 2280 5652 2286 5704
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5692 4675 5695
rect 4706 5692 4712 5704
rect 4663 5664 4712 5692
rect 4663 5661 4675 5664
rect 4617 5655 4675 5661
rect 2884 5556 2912 5655
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5692 8815 5695
rect 8846 5692 8852 5704
rect 8803 5664 8852 5692
rect 8803 5661 8815 5664
rect 8757 5655 8815 5661
rect 8846 5652 8852 5664
rect 8904 5652 8910 5704
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 4893 5627 4951 5633
rect 4893 5593 4905 5627
rect 4939 5624 4951 5627
rect 5718 5624 5724 5636
rect 4939 5596 5724 5624
rect 4939 5593 4951 5596
rect 4893 5587 4951 5593
rect 5718 5584 5724 5596
rect 5776 5584 5782 5636
rect 8110 5584 8116 5636
rect 8168 5624 8174 5636
rect 8956 5624 8984 5655
rect 8168 5596 8984 5624
rect 8168 5584 8174 5596
rect 3234 5556 3240 5568
rect 2884 5528 3240 5556
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 6730 5516 6736 5568
rect 6788 5556 6794 5568
rect 7745 5559 7803 5565
rect 7745 5556 7757 5559
rect 6788 5528 7757 5556
rect 6788 5516 6794 5528
rect 7745 5525 7757 5528
rect 7791 5525 7803 5559
rect 7745 5519 7803 5525
rect 8018 5516 8024 5568
rect 8076 5516 8082 5568
rect 8938 5516 8944 5568
rect 8996 5556 9002 5568
rect 9769 5559 9827 5565
rect 9769 5556 9781 5559
rect 8996 5528 9781 5556
rect 8996 5516 9002 5528
rect 9769 5525 9781 5528
rect 9815 5525 9827 5559
rect 9769 5519 9827 5525
rect 552 5466 10304 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 10304 5466
rect 552 5392 10304 5414
rect 6822 5352 6828 5364
rect 5920 5324 6828 5352
rect 1673 5287 1731 5293
rect 1673 5253 1685 5287
rect 1719 5284 1731 5287
rect 2222 5284 2228 5296
rect 1719 5256 2228 5284
rect 1719 5253 1731 5256
rect 1673 5247 1731 5253
rect 2222 5244 2228 5256
rect 2280 5284 2286 5296
rect 3418 5284 3424 5296
rect 2280 5256 3424 5284
rect 2280 5244 2286 5256
rect 3418 5244 3424 5256
rect 3476 5244 3482 5296
rect 4246 5244 4252 5296
rect 4304 5284 4310 5296
rect 4304 5256 4384 5284
rect 4304 5244 4310 5256
rect 4356 5225 4384 5256
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5216 4675 5219
rect 5810 5216 5816 5228
rect 4663 5188 5816 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 2777 5151 2835 5157
rect 2777 5117 2789 5151
rect 2823 5148 2835 5151
rect 3421 5151 3479 5157
rect 3421 5148 3433 5151
rect 2823 5120 3433 5148
rect 2823 5117 2835 5120
rect 2777 5111 2835 5117
rect 3421 5117 3433 5120
rect 3467 5148 3479 5151
rect 4246 5148 4252 5160
rect 3467 5120 4252 5148
rect 3467 5117 3479 5120
rect 3421 5111 3479 5117
rect 4246 5108 4252 5120
rect 4304 5108 4310 5160
rect 5718 5108 5724 5160
rect 5776 5108 5782 5160
rect 5920 5157 5948 5324
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7193 5355 7251 5361
rect 7193 5321 7205 5355
rect 7239 5352 7251 5355
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7239 5324 7389 5352
rect 7239 5321 7251 5324
rect 7193 5315 7251 5321
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 7377 5315 7435 5321
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 9953 5355 10011 5361
rect 9953 5352 9965 5355
rect 9916 5324 9965 5352
rect 9916 5312 9922 5324
rect 9953 5321 9965 5324
rect 9999 5321 10011 5355
rect 9953 5315 10011 5321
rect 6730 5284 6736 5296
rect 6012 5256 6736 5284
rect 6012 5157 6040 5256
rect 6730 5244 6736 5256
rect 6788 5244 6794 5296
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 6564 5188 8401 5216
rect 5905 5151 5963 5157
rect 5905 5117 5917 5151
rect 5951 5117 5963 5151
rect 5905 5111 5963 5117
rect 5997 5151 6055 5157
rect 5997 5117 6009 5151
rect 6043 5117 6055 5151
rect 5997 5111 6055 5117
rect 6086 5108 6092 5160
rect 6144 5108 6150 5160
rect 6564 5157 6592 5188
rect 8389 5185 8401 5188
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 8478 5176 8484 5228
rect 8536 5216 8542 5228
rect 8665 5219 8723 5225
rect 8665 5216 8677 5219
rect 8536 5188 8677 5216
rect 8536 5176 8542 5188
rect 8665 5185 8677 5188
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 8846 5176 8852 5228
rect 8904 5216 8910 5228
rect 9309 5219 9367 5225
rect 9309 5216 9321 5219
rect 8904 5188 9321 5216
rect 8904 5176 8910 5188
rect 9309 5185 9321 5188
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 6730 5157 6736 5160
rect 6273 5151 6331 5157
rect 6273 5117 6285 5151
rect 6319 5117 6331 5151
rect 6273 5111 6331 5117
rect 6549 5151 6607 5157
rect 6549 5117 6561 5151
rect 6595 5117 6607 5151
rect 6549 5111 6607 5117
rect 6697 5151 6736 5157
rect 6697 5117 6709 5151
rect 6697 5111 6736 5117
rect 1949 5083 2007 5089
rect 1949 5049 1961 5083
rect 1995 5080 2007 5083
rect 2133 5083 2191 5089
rect 2133 5080 2145 5083
rect 1995 5052 2145 5080
rect 1995 5049 2007 5052
rect 1949 5043 2007 5049
rect 2133 5049 2145 5052
rect 2179 5049 2191 5083
rect 2133 5043 2191 5049
rect 3142 5040 3148 5092
rect 3200 5080 3206 5092
rect 3237 5083 3295 5089
rect 3237 5080 3249 5083
rect 3200 5052 3249 5080
rect 3200 5040 3206 5052
rect 3237 5049 3249 5052
rect 3283 5080 3295 5083
rect 4522 5080 4528 5092
rect 3283 5052 4528 5080
rect 3283 5049 3295 5052
rect 3237 5043 3295 5049
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 1486 4972 1492 5024
rect 1544 4972 1550 5024
rect 3510 4972 3516 5024
rect 3568 5012 3574 5024
rect 3605 5015 3663 5021
rect 3605 5012 3617 5015
rect 3568 4984 3617 5012
rect 3568 4972 3574 4984
rect 3605 4981 3617 4984
rect 3651 4981 3663 5015
rect 3605 4975 3663 4981
rect 5350 4972 5356 5024
rect 5408 5012 5414 5024
rect 6288 5012 6316 5111
rect 6730 5108 6736 5111
rect 6788 5108 6794 5160
rect 7006 5108 7012 5160
rect 7064 5157 7070 5160
rect 7064 5148 7072 5157
rect 7064 5120 7109 5148
rect 7064 5111 7072 5120
rect 7064 5108 7070 5111
rect 7190 5108 7196 5160
rect 7248 5148 7254 5160
rect 7285 5151 7343 5157
rect 7285 5148 7297 5151
rect 7248 5120 7297 5148
rect 7248 5108 7254 5120
rect 7285 5117 7297 5120
rect 7331 5117 7343 5151
rect 7285 5111 7343 5117
rect 7653 5151 7711 5157
rect 7653 5117 7665 5151
rect 7699 5148 7711 5151
rect 7742 5148 7748 5160
rect 7699 5120 7748 5148
rect 7699 5117 7711 5120
rect 7653 5111 7711 5117
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 8202 5108 8208 5160
rect 8260 5148 8266 5160
rect 8757 5151 8815 5157
rect 8757 5148 8769 5151
rect 8260 5120 8769 5148
rect 8260 5108 8266 5120
rect 8757 5117 8769 5120
rect 8803 5117 8815 5151
rect 8757 5111 8815 5117
rect 6822 5040 6828 5092
rect 6880 5040 6886 5092
rect 6917 5083 6975 5089
rect 6917 5049 6929 5083
rect 6963 5049 6975 5083
rect 6917 5043 6975 5049
rect 5408 4984 6316 5012
rect 5408 4972 5414 4984
rect 6454 4972 6460 5024
rect 6512 4972 6518 5024
rect 6546 4972 6552 5024
rect 6604 5012 6610 5024
rect 6932 5012 6960 5043
rect 6604 4984 6960 5012
rect 7837 5015 7895 5021
rect 6604 4972 6610 4984
rect 7837 4981 7849 5015
rect 7883 5012 7895 5015
rect 8202 5012 8208 5024
rect 7883 4984 8208 5012
rect 7883 4981 7895 4984
rect 7837 4975 7895 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 552 4922 10304 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 10304 4922
rect 552 4848 10304 4870
rect 6914 4808 6920 4820
rect 6656 4780 6920 4808
rect 1204 4743 1262 4749
rect 1204 4709 1216 4743
rect 1250 4740 1262 4743
rect 1486 4740 1492 4752
rect 1250 4712 1492 4740
rect 1250 4709 1262 4712
rect 1204 4703 1262 4709
rect 1486 4700 1492 4712
rect 1544 4700 1550 4752
rect 4525 4743 4583 4749
rect 4525 4709 4537 4743
rect 4571 4740 4583 4743
rect 5534 4740 5540 4752
rect 4571 4712 5540 4740
rect 4571 4709 4583 4712
rect 4525 4703 4583 4709
rect 5534 4700 5540 4712
rect 5592 4700 5598 4752
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4641 2559 4675
rect 2501 4635 2559 4641
rect 2685 4675 2743 4681
rect 2685 4641 2697 4675
rect 2731 4672 2743 4675
rect 4154 4672 4160 4684
rect 2731 4644 4160 4672
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 934 4564 940 4616
rect 992 4564 998 4616
rect 2516 4604 2544 4635
rect 4154 4632 4160 4644
rect 4212 4632 4218 4684
rect 4430 4632 4436 4684
rect 4488 4672 4494 4684
rect 4617 4675 4675 4681
rect 4617 4672 4629 4675
rect 4488 4644 4629 4672
rect 4488 4632 4494 4644
rect 4617 4641 4629 4644
rect 4663 4641 4675 4675
rect 4617 4635 4675 4641
rect 4798 4632 4804 4684
rect 4856 4632 4862 4684
rect 5256 4675 5314 4681
rect 5256 4672 5268 4675
rect 5184 4644 5268 4672
rect 2774 4604 2780 4616
rect 2516 4576 2780 4604
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 952 4468 980 4564
rect 5184 4536 5212 4644
rect 5256 4641 5268 4644
rect 5302 4641 5314 4675
rect 5256 4635 5314 4641
rect 5350 4632 5356 4684
rect 5408 4632 5414 4684
rect 5442 4632 5448 4684
rect 5500 4632 5506 4684
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4641 5687 4675
rect 5629 4635 5687 4641
rect 6457 4675 6515 4681
rect 6457 4641 6469 4675
rect 6503 4672 6515 4675
rect 6546 4672 6552 4684
rect 6503 4644 6552 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 5644 4604 5672 4635
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 6656 4681 6684 4780
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 7466 4768 7472 4820
rect 7524 4768 7530 4820
rect 7742 4768 7748 4820
rect 7800 4768 7806 4820
rect 6730 4700 6736 4752
rect 6788 4740 6794 4752
rect 7484 4740 7512 4768
rect 8205 4743 8263 4749
rect 8205 4740 8217 4743
rect 6788 4712 7144 4740
rect 7484 4712 8217 4740
rect 6788 4700 6794 4712
rect 6641 4675 6699 4681
rect 6641 4641 6653 4675
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4674 6883 4675
rect 6914 4674 6920 4684
rect 6871 4646 6920 4674
rect 6871 4641 6883 4646
rect 6825 4635 6883 4641
rect 6914 4632 6920 4646
rect 6972 4632 6978 4684
rect 7116 4681 7144 4712
rect 8205 4709 8217 4712
rect 8251 4709 8263 4743
rect 8205 4703 8263 4709
rect 9766 4700 9772 4752
rect 9824 4700 9830 4752
rect 7282 4681 7288 4684
rect 7009 4675 7067 4681
rect 7009 4641 7021 4675
rect 7055 4641 7067 4675
rect 7009 4635 7067 4641
rect 7101 4675 7159 4681
rect 7101 4641 7113 4675
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 7249 4675 7288 4681
rect 7249 4641 7261 4675
rect 7249 4635 7288 4641
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 5644 4576 6745 4604
rect 6086 4536 6092 4548
rect 5184 4508 6092 4536
rect 6086 4496 6092 4508
rect 6144 4496 6150 4548
rect 1302 4468 1308 4480
rect 952 4440 1308 4468
rect 1302 4428 1308 4440
rect 1360 4428 1366 4480
rect 2314 4428 2320 4480
rect 2372 4428 2378 4480
rect 2593 4471 2651 4477
rect 2593 4437 2605 4471
rect 2639 4468 2651 4471
rect 3050 4468 3056 4480
rect 2639 4440 3056 4468
rect 2639 4437 2651 4440
rect 2593 4431 2651 4437
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 3234 4428 3240 4480
rect 3292 4428 3298 4480
rect 4706 4428 4712 4480
rect 4764 4428 4770 4480
rect 5626 4428 5632 4480
rect 5684 4428 5690 4480
rect 6270 4428 6276 4480
rect 6328 4428 6334 4480
rect 6564 4468 6592 4576
rect 6733 4573 6745 4576
rect 6779 4573 6791 4607
rect 7024 4604 7052 4635
rect 7282 4632 7288 4635
rect 7340 4632 7346 4684
rect 7374 4632 7380 4684
rect 7432 4632 7438 4684
rect 7466 4632 7472 4684
rect 7524 4632 7530 4684
rect 7558 4632 7564 4684
rect 7616 4681 7622 4684
rect 7616 4675 7665 4681
rect 7616 4641 7619 4675
rect 7653 4672 7665 4675
rect 8018 4672 8024 4684
rect 7653 4644 8024 4672
rect 7653 4641 7665 4644
rect 7616 4635 7665 4641
rect 7616 4632 7622 4635
rect 8018 4632 8024 4644
rect 8076 4632 8082 4684
rect 7834 4604 7840 4616
rect 7024 4576 7840 4604
rect 6733 4567 6791 4573
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 8018 4468 8024 4480
rect 6564 4440 8024 4468
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 552 4378 10304 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 10304 4378
rect 552 4304 10304 4326
rect 2685 4267 2743 4273
rect 2685 4233 2697 4267
rect 2731 4264 2743 4267
rect 3142 4264 3148 4276
rect 2731 4236 3148 4264
rect 2731 4233 2743 4236
rect 2685 4227 2743 4233
rect 3142 4224 3148 4236
rect 3200 4224 3206 4276
rect 3421 4267 3479 4273
rect 3421 4233 3433 4267
rect 3467 4264 3479 4267
rect 3510 4264 3516 4276
rect 3467 4236 3516 4264
rect 3467 4233 3479 4236
rect 3421 4227 3479 4233
rect 3510 4224 3516 4236
rect 3568 4224 3574 4276
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 4985 4267 5043 4273
rect 4985 4264 4997 4267
rect 4856 4236 4997 4264
rect 4856 4224 4862 4236
rect 4985 4233 4997 4236
rect 5031 4264 5043 4267
rect 6546 4264 6552 4276
rect 5031 4236 6552 4264
rect 5031 4233 5043 4236
rect 4985 4227 5043 4233
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 6917 4267 6975 4273
rect 6917 4233 6929 4267
rect 6963 4264 6975 4267
rect 7190 4264 7196 4276
rect 6963 4236 7196 4264
rect 6963 4233 6975 4236
rect 6917 4227 6975 4233
rect 7190 4224 7196 4236
rect 7248 4224 7254 4276
rect 7469 4267 7527 4273
rect 7469 4233 7481 4267
rect 7515 4264 7527 4267
rect 7558 4264 7564 4276
rect 7515 4236 7564 4264
rect 7515 4233 7527 4236
rect 7469 4227 7527 4233
rect 7558 4224 7564 4236
rect 7616 4224 7622 4276
rect 8481 4267 8539 4273
rect 8481 4233 8493 4267
rect 8527 4264 8539 4267
rect 8846 4264 8852 4276
rect 8527 4236 8852 4264
rect 8527 4233 8539 4236
rect 8481 4227 8539 4233
rect 8846 4224 8852 4236
rect 8904 4264 8910 4276
rect 9214 4264 9220 4276
rect 8904 4236 9220 4264
rect 8904 4224 8910 4236
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 2314 4156 2320 4208
rect 2372 4196 2378 4208
rect 4246 4196 4252 4208
rect 2372 4168 4252 4196
rect 2372 4156 2378 4168
rect 1302 4020 1308 4072
rect 1360 4020 1366 4072
rect 2700 4060 2728 4168
rect 4246 4156 4252 4168
rect 4304 4156 4310 4208
rect 6365 4199 6423 4205
rect 6365 4165 6377 4199
rect 6411 4196 6423 4199
rect 6454 4196 6460 4208
rect 6411 4168 6460 4196
rect 6411 4165 6423 4168
rect 6365 4159 6423 4165
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 2961 4131 3019 4137
rect 2961 4128 2973 4131
rect 2832 4100 2973 4128
rect 2832 4088 2838 4100
rect 2961 4097 2973 4100
rect 3007 4128 3019 4131
rect 4154 4128 4160 4140
rect 3007 4100 3740 4128
rect 3007 4097 3019 4100
rect 2961 4091 3019 4097
rect 2869 4063 2927 4069
rect 2869 4060 2881 4063
rect 2700 4032 2881 4060
rect 2869 4029 2881 4032
rect 2915 4029 2927 4063
rect 2869 4023 2927 4029
rect 3053 4063 3111 4069
rect 3053 4029 3065 4063
rect 3099 4060 3111 4063
rect 3142 4060 3148 4072
rect 3099 4032 3148 4060
rect 3099 4029 3111 4032
rect 3053 4023 3111 4029
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 3436 4001 3464 4100
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 3712 4069 3740 4100
rect 3896 4100 4160 4128
rect 3896 4069 3924 4100
rect 4154 4088 4160 4100
rect 4212 4128 4218 4140
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 4212 4100 5273 4128
rect 4212 4088 4218 4100
rect 5261 4097 5273 4100
rect 5307 4128 5319 4131
rect 5350 4128 5356 4140
rect 5307 4100 5356 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 7374 4128 7380 4140
rect 7208 4100 7380 4128
rect 3697 4063 3755 4069
rect 3568 4032 3648 4060
rect 3568 4020 3574 4032
rect 3620 4001 3648 4032
rect 3697 4029 3709 4063
rect 3743 4029 3755 4063
rect 3697 4023 3755 4029
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4029 3939 4063
rect 4430 4060 4436 4072
rect 3881 4023 3939 4029
rect 4080 4032 4436 4060
rect 1572 3995 1630 4001
rect 1572 3961 1584 3995
rect 1618 3992 1630 3995
rect 3405 3995 3464 4001
rect 1618 3964 3280 3992
rect 1618 3961 1630 3964
rect 1572 3955 1630 3961
rect 3252 3933 3280 3964
rect 3405 3961 3417 3995
rect 3451 3964 3464 3995
rect 3605 3995 3663 4001
rect 3451 3961 3463 3964
rect 3405 3955 3463 3961
rect 3605 3961 3617 3995
rect 3651 3961 3663 3995
rect 3605 3955 3663 3961
rect 3237 3927 3295 3933
rect 3237 3893 3249 3927
rect 3283 3893 3295 3927
rect 3237 3887 3295 3893
rect 3510 3884 3516 3936
rect 3568 3924 3574 3936
rect 4080 3933 4108 4032
rect 4430 4020 4436 4032
rect 4488 4020 4494 4072
rect 4617 4063 4675 4069
rect 4617 4029 4629 4063
rect 4663 4060 4675 4063
rect 5074 4060 5080 4072
rect 4663 4032 5080 4060
rect 4663 4029 4675 4032
rect 4617 4023 4675 4029
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 5169 4063 5227 4069
rect 5169 4029 5181 4063
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 4525 3995 4583 4001
rect 4525 3992 4537 3995
rect 4356 3964 4537 3992
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 3568 3896 4077 3924
rect 3568 3884 3574 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 4065 3887 4123 3893
rect 4154 3884 4160 3936
rect 4212 3924 4218 3936
rect 4356 3924 4384 3964
rect 4525 3961 4537 3964
rect 4571 3992 4583 3995
rect 5184 3992 5212 4023
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 7208 4069 7236 4100
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 6549 4063 6607 4069
rect 6549 4060 6561 4063
rect 6328 4032 6561 4060
rect 6328 4020 6334 4032
rect 6549 4029 6561 4032
rect 6595 4029 6607 4063
rect 6549 4023 6607 4029
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4029 7251 4063
rect 7193 4023 7251 4029
rect 7282 4020 7288 4072
rect 7340 4020 7346 4072
rect 7561 4063 7619 4069
rect 7561 4029 7573 4063
rect 7607 4029 7619 4063
rect 7561 4023 7619 4029
rect 4571 3964 5212 3992
rect 6641 3995 6699 4001
rect 4571 3961 4583 3964
rect 4525 3955 4583 3961
rect 6641 3961 6653 3995
rect 6687 3992 6699 3995
rect 7009 3995 7067 4001
rect 7009 3992 7021 3995
rect 6687 3964 7021 3992
rect 6687 3961 6699 3964
rect 6641 3955 6699 3961
rect 7009 3961 7021 3964
rect 7055 3961 7067 3995
rect 7009 3955 7067 3961
rect 7466 3952 7472 4004
rect 7524 3992 7530 4004
rect 7576 3992 7604 4023
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 9861 4063 9919 4069
rect 9861 4060 9873 4063
rect 9824 4032 9873 4060
rect 9824 4020 9830 4032
rect 9861 4029 9873 4032
rect 9907 4029 9919 4063
rect 9861 4023 9919 4029
rect 7524 3964 7604 3992
rect 7524 3952 7530 3964
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 9594 3995 9652 4001
rect 9594 3992 9606 3995
rect 9088 3964 9606 3992
rect 9088 3952 9094 3964
rect 9594 3961 9606 3964
rect 9640 3961 9652 3995
rect 9594 3955 9652 3961
rect 4212 3896 4384 3924
rect 4433 3927 4491 3933
rect 4212 3884 4218 3896
rect 4433 3893 4445 3927
rect 4479 3924 4491 3927
rect 4614 3924 4620 3936
rect 4479 3896 4620 3924
rect 4479 3893 4491 3896
rect 4433 3887 4491 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4798 3884 4804 3936
rect 4856 3884 4862 3936
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 6733 3927 6791 3933
rect 6733 3924 6745 3927
rect 5684 3896 6745 3924
rect 5684 3884 5690 3896
rect 6733 3893 6745 3896
rect 6779 3893 6791 3927
rect 6733 3887 6791 3893
rect 552 3834 10304 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 10304 3834
rect 552 3760 10304 3782
rect 3789 3723 3847 3729
rect 3789 3689 3801 3723
rect 3835 3720 3847 3723
rect 4154 3720 4160 3732
rect 3835 3692 4160 3720
rect 3835 3689 3847 3692
rect 3789 3683 3847 3689
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5261 3723 5319 3729
rect 5261 3720 5273 3723
rect 5132 3692 5273 3720
rect 5132 3680 5138 3692
rect 5261 3689 5273 3692
rect 5307 3689 5319 3723
rect 5261 3683 5319 3689
rect 7282 3680 7288 3732
rect 7340 3680 7346 3732
rect 7653 3723 7711 3729
rect 7653 3689 7665 3723
rect 7699 3720 7711 3723
rect 8662 3720 8668 3732
rect 7699 3692 8668 3720
rect 7699 3689 7711 3692
rect 7653 3683 7711 3689
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 9030 3680 9036 3732
rect 9088 3680 9094 3732
rect 1302 3612 1308 3664
rect 1360 3652 1366 3664
rect 3234 3652 3240 3664
rect 1360 3624 3240 3652
rect 1360 3612 1366 3624
rect 2424 3593 2452 3624
rect 3234 3612 3240 3624
rect 3292 3652 3298 3664
rect 3292 3624 3924 3652
rect 3292 3612 3298 3624
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3553 2467 3587
rect 2409 3547 2467 3553
rect 2676 3587 2734 3593
rect 2676 3553 2688 3587
rect 2722 3584 2734 3587
rect 3142 3584 3148 3596
rect 2722 3556 3148 3584
rect 2722 3553 2734 3556
rect 2676 3547 2734 3553
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 3896 3525 3924 3624
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 8938 3652 8944 3664
rect 8260 3624 8432 3652
rect 8260 3612 8266 3624
rect 4154 3593 4160 3596
rect 4148 3547 4160 3593
rect 4154 3544 4160 3547
rect 4212 3544 4218 3596
rect 7374 3544 7380 3596
rect 7432 3544 7438 3596
rect 7742 3544 7748 3596
rect 7800 3544 7806 3596
rect 7834 3544 7840 3596
rect 7892 3544 7898 3596
rect 8018 3544 8024 3596
rect 8076 3544 8082 3596
rect 8294 3544 8300 3596
rect 8352 3544 8358 3596
rect 8404 3593 8432 3624
rect 8792 3624 8944 3652
rect 8389 3587 8447 3593
rect 8389 3553 8401 3587
rect 8435 3553 8447 3587
rect 8389 3547 8447 3553
rect 8573 3587 8631 3593
rect 8573 3553 8585 3587
rect 8619 3553 8631 3587
rect 8573 3547 8631 3553
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3485 3939 3519
rect 3881 3479 3939 3485
rect 3896 3380 3924 3479
rect 7929 3451 7987 3457
rect 7929 3417 7941 3451
rect 7975 3448 7987 3451
rect 8386 3448 8392 3460
rect 7975 3420 8392 3448
rect 7975 3417 7987 3420
rect 7929 3411 7987 3417
rect 8386 3408 8392 3420
rect 8444 3408 8450 3460
rect 8588 3448 8616 3547
rect 8662 3544 8668 3596
rect 8720 3544 8726 3596
rect 8792 3593 8820 3624
rect 8938 3612 8944 3624
rect 8996 3612 9002 3664
rect 8792 3587 8861 3593
rect 8792 3556 8815 3587
rect 8803 3553 8815 3556
rect 8849 3553 8861 3587
rect 8803 3547 8861 3553
rect 9122 3544 9128 3596
rect 9180 3544 9186 3596
rect 9214 3544 9220 3596
rect 9272 3584 9278 3596
rect 9309 3587 9367 3593
rect 9309 3584 9321 3587
rect 9272 3556 9321 3584
rect 9272 3544 9278 3556
rect 9309 3553 9321 3556
rect 9355 3553 9367 3587
rect 9309 3547 9367 3553
rect 9493 3451 9551 3457
rect 9493 3448 9505 3451
rect 8588 3420 9505 3448
rect 9493 3417 9505 3420
rect 9539 3417 9551 3451
rect 9493 3411 9551 3417
rect 4246 3380 4252 3392
rect 3896 3352 4252 3380
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 8205 3383 8263 3389
rect 8205 3380 8217 3383
rect 8076 3352 8217 3380
rect 8076 3340 8082 3352
rect 8205 3349 8217 3352
rect 8251 3349 8263 3383
rect 8205 3343 8263 3349
rect 552 3290 10304 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 10304 3290
rect 552 3216 10304 3238
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 3237 3179 3295 3185
rect 3237 3176 3249 3179
rect 3200 3148 3249 3176
rect 3200 3136 3206 3148
rect 3237 3145 3249 3148
rect 3283 3145 3295 3179
rect 3237 3139 3295 3145
rect 3421 3179 3479 3185
rect 3421 3145 3433 3179
rect 3467 3176 3479 3179
rect 3510 3176 3516 3188
rect 3467 3148 3516 3176
rect 3467 3145 3479 3148
rect 3421 3139 3479 3145
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 3973 3179 4031 3185
rect 3973 3145 3985 3179
rect 4019 3176 4031 3179
rect 4062 3176 4068 3188
rect 4019 3148 4068 3176
rect 4019 3145 4031 3148
rect 3973 3139 4031 3145
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4157 3179 4215 3185
rect 4157 3145 4169 3179
rect 4203 3176 4215 3179
rect 4525 3179 4583 3185
rect 4525 3176 4537 3179
rect 4203 3148 4537 3176
rect 4203 3145 4215 3148
rect 4157 3139 4215 3145
rect 4525 3145 4537 3148
rect 4571 3145 4583 3179
rect 4525 3139 4583 3145
rect 8021 3179 8079 3185
rect 8021 3145 8033 3179
rect 8067 3176 8079 3179
rect 8294 3176 8300 3188
rect 8067 3148 8300 3176
rect 8067 3145 8079 3148
rect 8021 3139 8079 3145
rect 8294 3136 8300 3148
rect 8352 3176 8358 3188
rect 8481 3179 8539 3185
rect 8481 3176 8493 3179
rect 8352 3148 8493 3176
rect 8352 3136 8358 3148
rect 8481 3145 8493 3148
rect 8527 3145 8539 3179
rect 9122 3176 9128 3188
rect 8481 3139 8539 3145
rect 8588 3148 9128 3176
rect 7742 3068 7748 3120
rect 7800 3108 7806 3120
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 7800 3080 7849 3108
rect 7800 3068 7806 3080
rect 7837 3077 7849 3080
rect 7883 3108 7895 3111
rect 8588 3108 8616 3148
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 7883 3080 8616 3108
rect 7883 3077 7895 3080
rect 7837 3071 7895 3077
rect 8202 3040 8208 3052
rect 7668 3012 8208 3040
rect 4617 2975 4675 2981
rect 4617 2941 4629 2975
rect 4663 2972 4675 2975
rect 4798 2972 4804 2984
rect 4663 2944 4804 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 7668 2981 7696 3012
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 7653 2975 7711 2981
rect 7653 2941 7665 2975
rect 7699 2941 7711 2975
rect 7653 2935 7711 2941
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 9861 2975 9919 2981
rect 9861 2972 9873 2975
rect 9824 2944 9873 2972
rect 9824 2932 9830 2944
rect 9861 2941 9873 2944
rect 9907 2941 9919 2975
rect 9861 2935 9919 2941
rect 3050 2864 3056 2916
rect 3108 2904 3114 2916
rect 3389 2907 3447 2913
rect 3389 2904 3401 2907
rect 3108 2876 3401 2904
rect 3108 2864 3114 2876
rect 3389 2873 3401 2876
rect 3435 2873 3447 2907
rect 3389 2867 3447 2873
rect 3510 2864 3516 2916
rect 3568 2904 3574 2916
rect 3605 2907 3663 2913
rect 3605 2904 3617 2907
rect 3568 2876 3617 2904
rect 3568 2864 3574 2876
rect 3605 2873 3617 2876
rect 3651 2904 3663 2907
rect 4341 2907 4399 2913
rect 4341 2904 4353 2907
rect 3651 2876 4353 2904
rect 3651 2873 3663 2876
rect 3605 2867 3663 2873
rect 4341 2873 4353 2876
rect 4387 2904 4399 2907
rect 5626 2904 5632 2916
rect 4387 2876 5632 2904
rect 4387 2873 4399 2876
rect 4341 2867 4399 2873
rect 5626 2864 5632 2876
rect 5684 2904 5690 2916
rect 7282 2904 7288 2916
rect 5684 2876 7288 2904
rect 5684 2864 5690 2876
rect 7282 2864 7288 2876
rect 7340 2904 7346 2916
rect 7469 2907 7527 2913
rect 7469 2904 7481 2907
rect 7340 2876 7481 2904
rect 7340 2864 7346 2876
rect 7469 2873 7481 2876
rect 7515 2904 7527 2907
rect 8110 2904 8116 2916
rect 7515 2876 8116 2904
rect 7515 2873 7527 2876
rect 7469 2867 7527 2873
rect 8110 2864 8116 2876
rect 8168 2864 8174 2916
rect 8202 2864 8208 2916
rect 8260 2864 8266 2916
rect 8570 2864 8576 2916
rect 8628 2904 8634 2916
rect 9594 2907 9652 2913
rect 9594 2904 9606 2907
rect 8628 2876 9606 2904
rect 8628 2864 8634 2876
rect 9594 2873 9606 2876
rect 9640 2873 9652 2907
rect 9594 2867 9652 2873
rect 4141 2839 4199 2845
rect 4141 2805 4153 2839
rect 4187 2836 4199 2839
rect 4706 2836 4712 2848
rect 4187 2808 4712 2836
rect 4187 2805 4199 2808
rect 4141 2799 4199 2805
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 8018 2845 8024 2848
rect 8005 2839 8024 2845
rect 8005 2805 8017 2839
rect 8005 2799 8024 2805
rect 8018 2796 8024 2799
rect 8076 2796 8082 2848
rect 552 2746 10304 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 10304 2746
rect 552 2672 10304 2694
rect 6457 2635 6515 2641
rect 4908 2604 5948 2632
rect 4709 2499 4767 2505
rect 4709 2465 4721 2499
rect 4755 2465 4767 2499
rect 4709 2459 4767 2465
rect 4724 2428 4752 2459
rect 4798 2456 4804 2508
rect 4856 2496 4862 2508
rect 4908 2505 4936 2604
rect 5442 2573 5448 2576
rect 5429 2567 5448 2573
rect 5429 2533 5441 2567
rect 5429 2527 5448 2533
rect 5442 2524 5448 2527
rect 5500 2524 5506 2576
rect 5626 2524 5632 2576
rect 5684 2524 5690 2576
rect 5813 2567 5871 2573
rect 5813 2533 5825 2567
rect 5859 2533 5871 2567
rect 5920 2564 5948 2604
rect 6457 2601 6469 2635
rect 6503 2632 6515 2635
rect 6546 2632 6552 2644
rect 6503 2604 6552 2632
rect 6503 2601 6515 2604
rect 6457 2595 6515 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 7469 2635 7527 2641
rect 7469 2601 7481 2635
rect 7515 2632 7527 2635
rect 7834 2632 7840 2644
rect 7515 2604 7840 2632
rect 7515 2601 7527 2604
rect 7469 2595 7527 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 8570 2632 8576 2644
rect 8527 2604 8576 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 6013 2567 6071 2573
rect 6013 2564 6025 2567
rect 5920 2536 6025 2564
rect 5813 2527 5871 2533
rect 6013 2533 6025 2536
rect 6059 2564 6071 2567
rect 6641 2567 6699 2573
rect 6641 2564 6653 2567
rect 6059 2536 6653 2564
rect 6059 2533 6071 2536
rect 6013 2527 6071 2533
rect 6641 2533 6653 2536
rect 6687 2533 6699 2567
rect 7929 2567 7987 2573
rect 7929 2564 7941 2567
rect 6641 2527 6699 2533
rect 7300 2536 7941 2564
rect 4893 2499 4951 2505
rect 4893 2496 4905 2499
rect 4856 2468 4905 2496
rect 4856 2456 4862 2468
rect 4893 2465 4905 2468
rect 4939 2465 4951 2499
rect 4893 2459 4951 2465
rect 5828 2428 5856 2527
rect 7300 2505 7328 2536
rect 7929 2533 7941 2536
rect 7975 2564 7987 2567
rect 8018 2564 8024 2576
rect 7975 2536 8024 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 8018 2524 8024 2536
rect 8076 2524 8082 2576
rect 8110 2524 8116 2576
rect 8168 2524 8174 2576
rect 8329 2567 8387 2573
rect 8329 2533 8341 2567
rect 8375 2564 8387 2567
rect 8662 2564 8668 2576
rect 8375 2536 8668 2564
rect 8375 2533 8387 2536
rect 8329 2527 8387 2533
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2465 6607 2499
rect 6549 2459 6607 2465
rect 6825 2499 6883 2505
rect 6825 2465 6837 2499
rect 6871 2496 6883 2499
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 6871 2468 7205 2496
rect 6871 2465 6883 2468
rect 6825 2459 6883 2465
rect 7193 2465 7205 2468
rect 7239 2496 7251 2499
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 7239 2468 7297 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 6178 2428 6184 2440
rect 4724 2400 6184 2428
rect 6178 2388 6184 2400
rect 6236 2428 6242 2440
rect 6564 2428 6592 2459
rect 7374 2456 7380 2508
rect 7432 2496 7438 2508
rect 7469 2499 7527 2505
rect 7469 2496 7481 2499
rect 7432 2468 7481 2496
rect 7432 2456 7438 2468
rect 7469 2465 7481 2468
rect 7515 2496 7527 2499
rect 7745 2499 7803 2505
rect 7745 2496 7757 2499
rect 7515 2468 7757 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 7745 2465 7757 2468
rect 7791 2496 7803 2499
rect 8202 2496 8208 2508
rect 7791 2468 8208 2496
rect 7791 2465 7803 2468
rect 7745 2459 7803 2465
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 6638 2428 6644 2440
rect 6236 2400 6316 2428
rect 6564 2400 6644 2428
rect 6236 2388 6242 2400
rect 6288 2369 6316 2400
rect 6638 2388 6644 2400
rect 6696 2428 6702 2440
rect 8478 2428 8484 2440
rect 6696 2400 8484 2428
rect 6696 2388 6702 2400
rect 8478 2388 8484 2400
rect 8536 2388 8542 2440
rect 6273 2363 6331 2369
rect 6273 2329 6285 2363
rect 6319 2360 6331 2363
rect 7466 2360 7472 2372
rect 6319 2332 7472 2360
rect 6319 2329 6331 2332
rect 6273 2323 6331 2329
rect 7466 2320 7472 2332
rect 7524 2320 7530 2372
rect 4798 2252 4804 2304
rect 4856 2252 4862 2304
rect 5258 2252 5264 2304
rect 5316 2252 5322 2304
rect 5445 2295 5503 2301
rect 5445 2261 5457 2295
rect 5491 2292 5503 2295
rect 5902 2292 5908 2304
rect 5491 2264 5908 2292
rect 5491 2261 5503 2264
rect 5445 2255 5503 2261
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 5994 2252 6000 2304
rect 6052 2252 6058 2304
rect 6181 2295 6239 2301
rect 6181 2261 6193 2295
rect 6227 2292 6239 2295
rect 6454 2292 6460 2304
rect 6227 2264 6460 2292
rect 6227 2261 6239 2264
rect 6181 2255 6239 2261
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 7098 2252 7104 2304
rect 7156 2252 7162 2304
rect 7561 2295 7619 2301
rect 7561 2261 7573 2295
rect 7607 2292 7619 2295
rect 7742 2292 7748 2304
rect 7607 2264 7748 2292
rect 7607 2261 7619 2264
rect 7561 2255 7619 2261
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 8297 2295 8355 2301
rect 8297 2261 8309 2295
rect 8343 2292 8355 2295
rect 8386 2292 8392 2304
rect 8343 2264 8392 2292
rect 8343 2261 8355 2264
rect 8297 2255 8355 2261
rect 8386 2252 8392 2264
rect 8444 2252 8450 2304
rect 552 2202 10304 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 10304 2202
rect 552 2128 10304 2150
rect 4249 2091 4307 2097
rect 4249 2057 4261 2091
rect 4295 2088 4307 2091
rect 4798 2088 4804 2100
rect 4295 2060 4804 2088
rect 4295 2057 4307 2060
rect 4249 2051 4307 2057
rect 4798 2048 4804 2060
rect 4856 2048 4862 2100
rect 5994 2048 6000 2100
rect 6052 2088 6058 2100
rect 6365 2091 6423 2097
rect 6365 2088 6377 2091
rect 6052 2060 6377 2088
rect 6052 2048 6058 2060
rect 6365 2057 6377 2060
rect 6411 2088 6423 2091
rect 6546 2088 6552 2100
rect 6411 2060 6552 2088
rect 6411 2057 6423 2060
rect 6365 2051 6423 2057
rect 6546 2048 6552 2060
rect 6604 2048 6610 2100
rect 6825 2091 6883 2097
rect 6825 2057 6837 2091
rect 6871 2088 6883 2091
rect 7101 2091 7159 2097
rect 7101 2088 7113 2091
rect 6871 2060 7113 2088
rect 6871 2057 6883 2060
rect 6825 2051 6883 2057
rect 7101 2057 7113 2060
rect 7147 2057 7159 2091
rect 7101 2051 7159 2057
rect 7742 2048 7748 2100
rect 7800 2048 7806 2100
rect 8202 2048 8208 2100
rect 8260 2088 8266 2100
rect 8389 2091 8447 2097
rect 8389 2088 8401 2091
rect 8260 2060 8401 2088
rect 8260 2048 8266 2060
rect 8389 2057 8401 2060
rect 8435 2057 8447 2091
rect 8389 2051 8447 2057
rect 4246 1912 4252 1964
rect 4304 1952 4310 1964
rect 4985 1955 5043 1961
rect 4985 1952 4997 1955
rect 4304 1924 4997 1952
rect 4304 1912 4310 1924
rect 4985 1921 4997 1924
rect 5031 1921 5043 1955
rect 4985 1915 5043 1921
rect 4890 1844 4896 1896
rect 4948 1844 4954 1896
rect 5258 1893 5264 1896
rect 5252 1884 5264 1893
rect 5219 1856 5264 1884
rect 5252 1847 5264 1856
rect 5258 1844 5264 1847
rect 5316 1844 5322 1896
rect 6454 1844 6460 1896
rect 6512 1844 6518 1896
rect 6638 1844 6644 1896
rect 6696 1844 6702 1896
rect 9766 1844 9772 1896
rect 9824 1844 9830 1896
rect 3510 1776 3516 1828
rect 3568 1816 3574 1828
rect 4065 1819 4123 1825
rect 4065 1816 4077 1819
rect 3568 1788 4077 1816
rect 3568 1776 3574 1788
rect 4065 1785 4077 1788
rect 4111 1785 4123 1819
rect 4065 1779 4123 1785
rect 4281 1819 4339 1825
rect 4281 1785 4293 1819
rect 4327 1816 4339 1819
rect 4525 1819 4583 1825
rect 4525 1816 4537 1819
rect 4327 1788 4537 1816
rect 4327 1785 4339 1788
rect 4281 1779 4339 1785
rect 4525 1785 4537 1788
rect 4571 1785 4583 1819
rect 4525 1779 4583 1785
rect 4709 1819 4767 1825
rect 4709 1785 4721 1819
rect 4755 1816 4767 1819
rect 6178 1816 6184 1828
rect 4755 1788 6184 1816
rect 4755 1785 4767 1788
rect 4709 1779 4767 1785
rect 6178 1776 6184 1788
rect 6236 1776 6242 1828
rect 7098 1825 7104 1828
rect 7085 1819 7104 1825
rect 7085 1785 7097 1819
rect 7085 1779 7104 1785
rect 7098 1776 7104 1779
rect 7156 1776 7162 1828
rect 7282 1776 7288 1828
rect 7340 1816 7346 1828
rect 7834 1825 7840 1828
rect 7561 1819 7619 1825
rect 7561 1816 7573 1819
rect 7340 1788 7573 1816
rect 7340 1776 7346 1788
rect 7561 1785 7573 1788
rect 7607 1785 7619 1819
rect 7561 1779 7619 1785
rect 7777 1819 7840 1825
rect 7777 1785 7789 1819
rect 7823 1785 7840 1819
rect 7777 1779 7840 1785
rect 7834 1776 7840 1779
rect 7892 1776 7898 1828
rect 9502 1819 9560 1825
rect 9502 1816 9514 1819
rect 7944 1788 9514 1816
rect 4154 1708 4160 1760
rect 4212 1748 4218 1760
rect 4433 1751 4491 1757
rect 4433 1748 4445 1751
rect 4212 1720 4445 1748
rect 4212 1708 4218 1720
rect 4433 1717 4445 1720
rect 4479 1717 4491 1751
rect 4433 1711 4491 1717
rect 6914 1708 6920 1760
rect 6972 1708 6978 1760
rect 7944 1757 7972 1788
rect 9502 1785 9514 1788
rect 9548 1785 9560 1819
rect 9502 1779 9560 1785
rect 7929 1751 7987 1757
rect 7929 1717 7941 1751
rect 7975 1717 7987 1751
rect 7929 1711 7987 1717
rect 552 1658 10304 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 10304 1658
rect 552 1584 10304 1606
rect 5902 1504 5908 1556
rect 5960 1544 5966 1556
rect 6457 1547 6515 1553
rect 6457 1544 6469 1547
rect 5960 1516 6469 1544
rect 5960 1504 5966 1516
rect 6457 1513 6469 1516
rect 6503 1513 6515 1547
rect 6457 1507 6515 1513
rect 6638 1504 6644 1556
rect 6696 1544 6702 1556
rect 6825 1547 6883 1553
rect 6825 1544 6837 1547
rect 6696 1516 6837 1544
rect 6696 1504 6702 1516
rect 6825 1513 6837 1516
rect 6871 1513 6883 1547
rect 6825 1507 6883 1513
rect 4154 1436 4160 1488
rect 4212 1476 4218 1488
rect 4505 1479 4563 1485
rect 4505 1476 4517 1479
rect 4212 1448 4517 1476
rect 4212 1436 4218 1448
rect 4505 1445 4517 1448
rect 4551 1445 4563 1479
rect 4505 1439 4563 1445
rect 4890 1436 4896 1488
rect 4948 1476 4954 1488
rect 4948 1448 6316 1476
rect 4948 1436 4954 1448
rect 4246 1368 4252 1420
rect 4304 1368 4310 1420
rect 5994 1368 6000 1420
rect 6052 1368 6058 1420
rect 6178 1408 6184 1420
rect 6104 1380 6184 1408
rect 5442 1300 5448 1352
rect 5500 1340 5506 1352
rect 5813 1343 5871 1349
rect 5813 1340 5825 1343
rect 5500 1312 5825 1340
rect 5500 1300 5506 1312
rect 5813 1309 5825 1312
rect 5859 1309 5871 1343
rect 5813 1303 5871 1309
rect 5629 1275 5687 1281
rect 5629 1241 5641 1275
rect 5675 1272 5687 1275
rect 6104 1272 6132 1380
rect 6178 1368 6184 1380
rect 6236 1368 6242 1420
rect 6288 1417 6316 1448
rect 6914 1436 6920 1488
rect 6972 1476 6978 1488
rect 7938 1479 7996 1485
rect 7938 1476 7950 1479
rect 6972 1448 7950 1476
rect 6972 1436 6978 1448
rect 7938 1445 7950 1448
rect 7984 1445 7996 1479
rect 7938 1439 7996 1445
rect 6273 1411 6331 1417
rect 6273 1377 6285 1411
rect 6319 1377 6331 1411
rect 6273 1371 6331 1377
rect 6365 1411 6423 1417
rect 6365 1377 6377 1411
rect 6411 1408 6423 1411
rect 6454 1408 6460 1420
rect 6411 1380 6460 1408
rect 6411 1377 6423 1380
rect 6365 1371 6423 1377
rect 6454 1368 6460 1380
rect 6512 1368 6518 1420
rect 8205 1343 8263 1349
rect 8205 1309 8217 1343
rect 8251 1340 8263 1343
rect 9766 1340 9772 1352
rect 8251 1312 9772 1340
rect 8251 1309 8263 1312
rect 8205 1303 8263 1309
rect 9766 1300 9772 1312
rect 9824 1300 9830 1352
rect 5675 1244 6132 1272
rect 5675 1241 5687 1244
rect 5629 1235 5687 1241
rect 552 1114 10304 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 10304 1114
rect 552 1040 10304 1062
rect 2682 892 2688 944
rect 2740 932 2746 944
rect 2777 935 2835 941
rect 2777 932 2789 935
rect 2740 904 2789 932
rect 2740 892 2746 904
rect 2777 901 2789 904
rect 2823 901 2835 935
rect 2777 895 2835 901
rect 8110 892 8116 944
rect 8168 932 8174 944
rect 8573 935 8631 941
rect 8573 932 8585 935
rect 8168 904 8585 932
rect 8168 892 8174 904
rect 8573 901 8585 904
rect 8619 901 8631 935
rect 8573 895 8631 901
rect 2958 756 2964 808
rect 3016 756 3022 808
rect 7650 756 7656 808
rect 7708 796 7714 808
rect 8389 799 8447 805
rect 8389 796 8401 799
rect 7708 768 8401 796
rect 7708 756 7714 768
rect 8389 765 8401 768
rect 8435 765 8447 799
rect 8389 759 8447 765
rect 552 570 10304 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 10304 570
rect 552 496 10304 518
<< via1 >>
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 2964 9460 3016 9512
rect 3516 9460 3568 9512
rect 4528 9664 4580 9716
rect 4160 9503 4212 9512
rect 4160 9469 4169 9503
rect 4169 9469 4203 9503
rect 4203 9469 4212 9503
rect 4160 9460 4212 9469
rect 5632 9460 5684 9512
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 9956 9460 10008 9512
rect 1124 9435 1176 9444
rect 1124 9401 1158 9435
rect 1158 9401 1176 9435
rect 1124 9392 1176 9401
rect 1216 9392 1268 9444
rect 2320 9367 2372 9376
rect 2320 9333 2329 9367
rect 2329 9333 2363 9367
rect 2363 9333 2372 9367
rect 2320 9324 2372 9333
rect 3240 9367 3292 9376
rect 3240 9333 3249 9367
rect 3249 9333 3283 9367
rect 3283 9333 3292 9367
rect 3240 9324 3292 9333
rect 3516 9324 3568 9376
rect 7748 9392 7800 9444
rect 5816 9324 5868 9376
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 7380 9324 7432 9376
rect 8116 9324 8168 9376
rect 8484 9392 8536 9444
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 1032 9027 1084 9036
rect 1032 8993 1041 9027
rect 1041 8993 1075 9027
rect 1075 8993 1084 9027
rect 1032 8984 1084 8993
rect 5632 9163 5684 9172
rect 5632 9129 5641 9163
rect 5641 9129 5675 9163
rect 5675 9129 5684 9163
rect 5632 9120 5684 9129
rect 3240 9052 3292 9104
rect 1216 8916 1268 8968
rect 5724 8984 5776 9036
rect 6828 9052 6880 9104
rect 6736 8984 6788 9036
rect 7012 8984 7064 9036
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 8668 8984 8720 9036
rect 4160 8916 4212 8968
rect 9956 8916 10008 8968
rect 2688 8823 2740 8832
rect 2688 8789 2697 8823
rect 2697 8789 2731 8823
rect 2731 8789 2740 8823
rect 2688 8780 2740 8789
rect 4252 8780 4304 8832
rect 7288 8823 7340 8832
rect 7288 8789 7297 8823
rect 7297 8789 7331 8823
rect 7331 8789 7340 8823
rect 7288 8780 7340 8789
rect 7656 8780 7708 8832
rect 9404 8780 9456 8832
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 1124 8576 1176 8628
rect 5724 8576 5776 8628
rect 6736 8576 6788 8628
rect 7748 8576 7800 8628
rect 5632 8508 5684 8560
rect 1216 8440 1268 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 6184 8440 6236 8492
rect 388 8372 440 8424
rect 5080 8415 5132 8424
rect 5080 8381 5089 8415
rect 5089 8381 5123 8415
rect 5123 8381 5132 8415
rect 5080 8372 5132 8381
rect 5356 8372 5408 8424
rect 7288 8440 7340 8492
rect 7932 8372 7984 8424
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 2044 8304 2096 8356
rect 5540 8304 5592 8356
rect 7840 8304 7892 8356
rect 9680 8347 9732 8356
rect 9680 8313 9698 8347
rect 9698 8313 9732 8347
rect 9680 8304 9732 8313
rect 3056 8279 3108 8288
rect 3056 8245 3065 8279
rect 3065 8245 3099 8279
rect 3099 8245 3108 8279
rect 3056 8236 3108 8245
rect 4160 8236 4212 8288
rect 5724 8279 5776 8288
rect 5724 8245 5733 8279
rect 5733 8245 5767 8279
rect 5767 8245 5776 8279
rect 5724 8236 5776 8245
rect 6460 8279 6512 8288
rect 6460 8245 6469 8279
rect 6469 8245 6503 8279
rect 6503 8245 6512 8279
rect 6460 8236 6512 8245
rect 7104 8236 7156 8288
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 5080 8032 5132 8084
rect 9680 8032 9732 8084
rect 2320 7964 2372 8016
rect 3516 7964 3568 8016
rect 1216 7896 1268 7948
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 4160 7896 4212 7948
rect 5632 7939 5684 7948
rect 5632 7905 5641 7939
rect 5641 7905 5675 7939
rect 5675 7905 5684 7939
rect 5632 7896 5684 7905
rect 6552 7896 6604 7948
rect 6828 7896 6880 7948
rect 7656 7939 7708 7948
rect 7656 7905 7690 7939
rect 7690 7905 7708 7939
rect 7656 7896 7708 7905
rect 9496 7896 9548 7948
rect 8392 7828 8444 7880
rect 2780 7692 2832 7744
rect 3332 7735 3384 7744
rect 3332 7701 3341 7735
rect 3341 7701 3375 7735
rect 3375 7701 3384 7735
rect 3332 7692 3384 7701
rect 4988 7735 5040 7744
rect 4988 7701 4997 7735
rect 4997 7701 5031 7735
rect 5031 7701 5040 7735
rect 4988 7692 5040 7701
rect 7288 7692 7340 7744
rect 8024 7692 8076 7744
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 8392 7531 8444 7540
rect 8392 7497 8401 7531
rect 8401 7497 8435 7531
rect 8435 7497 8444 7531
rect 8392 7488 8444 7497
rect 2780 7395 2832 7404
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 2780 7352 2832 7361
rect 3056 7352 3108 7404
rect 4252 7420 4304 7472
rect 6828 7395 6880 7404
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 2044 7327 2096 7336
rect 2044 7293 2053 7327
rect 2053 7293 2087 7327
rect 2087 7293 2096 7327
rect 2044 7284 2096 7293
rect 2504 7284 2556 7336
rect 4252 7284 4304 7336
rect 5724 7284 5776 7336
rect 7104 7327 7156 7336
rect 7104 7293 7138 7327
rect 7138 7293 7156 7327
rect 7104 7284 7156 7293
rect 9772 7327 9824 7336
rect 9772 7293 9781 7327
rect 9781 7293 9815 7327
rect 9815 7293 9824 7327
rect 9772 7284 9824 7293
rect 9404 7216 9456 7268
rect 1308 7148 1360 7200
rect 2412 7191 2464 7200
rect 2412 7157 2421 7191
rect 2421 7157 2455 7191
rect 2455 7157 2464 7191
rect 2412 7148 2464 7157
rect 3516 7148 3568 7200
rect 4804 7191 4856 7200
rect 4804 7157 4813 7191
rect 4813 7157 4847 7191
rect 4847 7157 4856 7191
rect 4804 7148 4856 7157
rect 7012 7148 7064 7200
rect 8208 7191 8260 7200
rect 8208 7157 8217 7191
rect 8217 7157 8251 7191
rect 8251 7157 8260 7191
rect 8208 7148 8260 7157
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 1216 6851 1268 6860
rect 1216 6817 1225 6851
rect 1225 6817 1259 6851
rect 1259 6817 1268 6851
rect 1216 6808 1268 6817
rect 2504 6740 2556 6792
rect 3424 6808 3476 6860
rect 4804 6876 4856 6928
rect 4160 6851 4212 6860
rect 4160 6817 4169 6851
rect 4169 6817 4203 6851
rect 4203 6817 4212 6851
rect 4160 6808 4212 6817
rect 4988 6808 5040 6860
rect 6828 6876 6880 6928
rect 9496 6876 9548 6928
rect 6460 6808 6512 6860
rect 8024 6808 8076 6860
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 9956 6851 10008 6860
rect 9956 6817 9965 6851
rect 9965 6817 9999 6851
rect 9999 6817 10008 6851
rect 9956 6808 10008 6817
rect 2964 6604 3016 6656
rect 3056 6604 3108 6656
rect 6092 6604 6144 6656
rect 7104 6604 7156 6656
rect 7932 6604 7984 6656
rect 8668 6604 8720 6656
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 3424 6400 3476 6452
rect 7932 6400 7984 6452
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 4712 6264 4764 6316
rect 7012 6307 7064 6316
rect 7012 6273 7021 6307
rect 7021 6273 7055 6307
rect 7055 6273 7064 6307
rect 7012 6264 7064 6273
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 7656 6264 7708 6316
rect 9772 6307 9824 6316
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 940 6239 992 6248
rect 940 6205 949 6239
rect 949 6205 983 6239
rect 983 6205 992 6239
rect 940 6196 992 6205
rect 3240 6239 3292 6248
rect 3240 6205 3249 6239
rect 3249 6205 3283 6239
rect 3283 6205 3292 6239
rect 3240 6196 3292 6205
rect 3516 6239 3568 6248
rect 3516 6205 3550 6239
rect 3550 6205 3568 6239
rect 3516 6196 3568 6205
rect 4252 6196 4304 6248
rect 7104 6239 7156 6248
rect 7104 6205 7138 6239
rect 7138 6205 7156 6239
rect 7104 6196 7156 6205
rect 1308 6128 1360 6180
rect 9496 6171 9548 6180
rect 9496 6137 9514 6171
rect 9514 6137 9548 6171
rect 9496 6128 9548 6137
rect 7104 6060 7156 6112
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 2044 5856 2096 5908
rect 2412 5856 2464 5908
rect 3056 5856 3108 5908
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 7840 5856 7892 5908
rect 9496 5856 9548 5908
rect 3332 5788 3384 5840
rect 5540 5788 5592 5840
rect 7472 5788 7524 5840
rect 10324 5788 10376 5840
rect 4528 5763 4580 5772
rect 4528 5729 4537 5763
rect 4537 5729 4571 5763
rect 4571 5729 4580 5763
rect 4528 5720 4580 5729
rect 7288 5720 7340 5772
rect 7932 5763 7984 5772
rect 7932 5729 7941 5763
rect 7941 5729 7975 5763
rect 7975 5729 7984 5763
rect 7932 5720 7984 5729
rect 8668 5763 8720 5772
rect 8668 5729 8677 5763
rect 8677 5729 8711 5763
rect 8711 5729 8720 5763
rect 8668 5720 8720 5729
rect 9864 5763 9916 5772
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 9864 5720 9916 5729
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 4712 5652 4764 5704
rect 8852 5652 8904 5704
rect 5724 5584 5776 5636
rect 8116 5584 8168 5636
rect 3240 5516 3292 5568
rect 6736 5516 6788 5568
rect 8024 5559 8076 5568
rect 8024 5525 8033 5559
rect 8033 5525 8067 5559
rect 8067 5525 8076 5559
rect 8024 5516 8076 5525
rect 8944 5516 8996 5568
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 2228 5244 2280 5296
rect 3424 5244 3476 5296
rect 4252 5244 4304 5296
rect 5816 5176 5868 5228
rect 4252 5151 4304 5160
rect 4252 5117 4261 5151
rect 4261 5117 4295 5151
rect 4295 5117 4304 5151
rect 4252 5108 4304 5117
rect 5724 5151 5776 5160
rect 5724 5117 5733 5151
rect 5733 5117 5767 5151
rect 5767 5117 5776 5151
rect 5724 5108 5776 5117
rect 6828 5312 6880 5364
rect 9864 5312 9916 5364
rect 6736 5244 6788 5296
rect 6092 5151 6144 5160
rect 6092 5117 6101 5151
rect 6101 5117 6135 5151
rect 6135 5117 6144 5151
rect 6092 5108 6144 5117
rect 8484 5176 8536 5228
rect 8852 5176 8904 5228
rect 6736 5151 6788 5160
rect 6736 5117 6743 5151
rect 6743 5117 6788 5151
rect 3148 5040 3200 5092
rect 4528 5040 4580 5092
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 3516 4972 3568 5024
rect 5356 4972 5408 5024
rect 6736 5108 6788 5117
rect 7012 5151 7064 5160
rect 7012 5117 7026 5151
rect 7026 5117 7060 5151
rect 7060 5117 7064 5151
rect 7012 5108 7064 5117
rect 7196 5108 7248 5160
rect 7748 5108 7800 5160
rect 8208 5108 8260 5160
rect 6828 5083 6880 5092
rect 6828 5049 6837 5083
rect 6837 5049 6871 5083
rect 6871 5049 6880 5083
rect 6828 5040 6880 5049
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 6552 4972 6604 5024
rect 8208 4972 8260 5024
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 1492 4700 1544 4752
rect 5540 4700 5592 4752
rect 940 4607 992 4616
rect 940 4573 949 4607
rect 949 4573 983 4607
rect 983 4573 992 4607
rect 940 4564 992 4573
rect 4160 4632 4212 4684
rect 4436 4632 4488 4684
rect 4804 4675 4856 4684
rect 4804 4641 4813 4675
rect 4813 4641 4847 4675
rect 4847 4641 4856 4675
rect 4804 4632 4856 4641
rect 2780 4564 2832 4616
rect 5356 4675 5408 4684
rect 5356 4641 5365 4675
rect 5365 4641 5399 4675
rect 5399 4641 5408 4675
rect 5356 4632 5408 4641
rect 5448 4675 5500 4684
rect 5448 4641 5457 4675
rect 5457 4641 5491 4675
rect 5491 4641 5500 4675
rect 5448 4632 5500 4641
rect 6552 4632 6604 4684
rect 6920 4768 6972 4820
rect 7472 4768 7524 4820
rect 7748 4811 7800 4820
rect 7748 4777 7757 4811
rect 7757 4777 7791 4811
rect 7791 4777 7800 4811
rect 7748 4768 7800 4777
rect 6736 4700 6788 4752
rect 6920 4632 6972 4684
rect 9772 4743 9824 4752
rect 9772 4709 9781 4743
rect 9781 4709 9815 4743
rect 9815 4709 9824 4743
rect 9772 4700 9824 4709
rect 7288 4675 7340 4684
rect 7288 4641 7295 4675
rect 7295 4641 7340 4675
rect 6092 4496 6144 4548
rect 1308 4428 1360 4480
rect 2320 4471 2372 4480
rect 2320 4437 2329 4471
rect 2329 4437 2363 4471
rect 2363 4437 2372 4471
rect 2320 4428 2372 4437
rect 3056 4428 3108 4480
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 4712 4471 4764 4480
rect 4712 4437 4721 4471
rect 4721 4437 4755 4471
rect 4755 4437 4764 4471
rect 4712 4428 4764 4437
rect 5632 4471 5684 4480
rect 5632 4437 5641 4471
rect 5641 4437 5675 4471
rect 5675 4437 5684 4471
rect 5632 4428 5684 4437
rect 6276 4471 6328 4480
rect 6276 4437 6285 4471
rect 6285 4437 6319 4471
rect 6319 4437 6328 4471
rect 6276 4428 6328 4437
rect 7288 4632 7340 4641
rect 7380 4675 7432 4684
rect 7380 4641 7389 4675
rect 7389 4641 7423 4675
rect 7423 4641 7432 4675
rect 7380 4632 7432 4641
rect 7472 4675 7524 4684
rect 7472 4641 7481 4675
rect 7481 4641 7515 4675
rect 7515 4641 7524 4675
rect 7472 4632 7524 4641
rect 7564 4632 7616 4684
rect 8024 4632 8076 4684
rect 7840 4564 7892 4616
rect 8024 4428 8076 4480
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 3148 4224 3200 4276
rect 3516 4224 3568 4276
rect 4804 4224 4856 4276
rect 6552 4224 6604 4276
rect 7196 4224 7248 4276
rect 7564 4224 7616 4276
rect 8852 4224 8904 4276
rect 9220 4224 9272 4276
rect 2320 4156 2372 4208
rect 4252 4199 4304 4208
rect 1308 4063 1360 4072
rect 1308 4029 1317 4063
rect 1317 4029 1351 4063
rect 1351 4029 1360 4063
rect 1308 4020 1360 4029
rect 4252 4165 4261 4199
rect 4261 4165 4295 4199
rect 4295 4165 4304 4199
rect 4252 4156 4304 4165
rect 6460 4156 6512 4208
rect 2780 4088 2832 4140
rect 3148 4020 3200 4072
rect 3516 4020 3568 4072
rect 4160 4088 4212 4140
rect 5356 4088 5408 4140
rect 3516 3884 3568 3936
rect 4436 4020 4488 4072
rect 5080 4063 5132 4072
rect 5080 4029 5089 4063
rect 5089 4029 5123 4063
rect 5123 4029 5132 4063
rect 5080 4020 5132 4029
rect 4160 3884 4212 3936
rect 6276 4020 6328 4072
rect 7380 4088 7432 4140
rect 7288 4063 7340 4072
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 7472 3952 7524 4004
rect 9772 4020 9824 4072
rect 9036 3952 9088 4004
rect 4620 3884 4672 3936
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 5632 3884 5684 3936
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 4160 3680 4212 3732
rect 5080 3680 5132 3732
rect 7288 3723 7340 3732
rect 7288 3689 7297 3723
rect 7297 3689 7331 3723
rect 7331 3689 7340 3723
rect 7288 3680 7340 3689
rect 8668 3680 8720 3732
rect 9036 3723 9088 3732
rect 9036 3689 9045 3723
rect 9045 3689 9079 3723
rect 9079 3689 9088 3723
rect 9036 3680 9088 3689
rect 1308 3612 1360 3664
rect 3240 3612 3292 3664
rect 3148 3544 3200 3596
rect 8208 3612 8260 3664
rect 4160 3587 4212 3596
rect 4160 3553 4194 3587
rect 4194 3553 4212 3587
rect 4160 3544 4212 3553
rect 7380 3587 7432 3596
rect 7380 3553 7389 3587
rect 7389 3553 7423 3587
rect 7423 3553 7432 3587
rect 7380 3544 7432 3553
rect 7748 3587 7800 3596
rect 7748 3553 7757 3587
rect 7757 3553 7791 3587
rect 7791 3553 7800 3587
rect 7748 3544 7800 3553
rect 7840 3587 7892 3596
rect 7840 3553 7849 3587
rect 7849 3553 7883 3587
rect 7883 3553 7892 3587
rect 7840 3544 7892 3553
rect 8024 3587 8076 3596
rect 8024 3553 8033 3587
rect 8033 3553 8067 3587
rect 8067 3553 8076 3587
rect 8024 3544 8076 3553
rect 8300 3587 8352 3596
rect 8300 3553 8309 3587
rect 8309 3553 8343 3587
rect 8343 3553 8352 3587
rect 8300 3544 8352 3553
rect 8392 3408 8444 3460
rect 8668 3587 8720 3596
rect 8668 3553 8677 3587
rect 8677 3553 8711 3587
rect 8711 3553 8720 3587
rect 8668 3544 8720 3553
rect 8944 3612 8996 3664
rect 9128 3587 9180 3596
rect 9128 3553 9137 3587
rect 9137 3553 9171 3587
rect 9171 3553 9180 3587
rect 9128 3544 9180 3553
rect 9220 3544 9272 3596
rect 4252 3340 4304 3392
rect 8024 3340 8076 3392
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 3148 3136 3200 3188
rect 3516 3136 3568 3188
rect 4068 3136 4120 3188
rect 8300 3136 8352 3188
rect 7748 3068 7800 3120
rect 9128 3136 9180 3188
rect 4804 2932 4856 2984
rect 8208 3000 8260 3052
rect 9772 2932 9824 2984
rect 3056 2864 3108 2916
rect 3516 2864 3568 2916
rect 5632 2864 5684 2916
rect 7288 2864 7340 2916
rect 8116 2864 8168 2916
rect 8208 2907 8260 2916
rect 8208 2873 8217 2907
rect 8217 2873 8251 2907
rect 8251 2873 8260 2907
rect 8208 2864 8260 2873
rect 8576 2864 8628 2916
rect 4712 2796 4764 2848
rect 8024 2839 8076 2848
rect 8024 2805 8051 2839
rect 8051 2805 8076 2839
rect 8024 2796 8076 2805
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 4804 2456 4856 2508
rect 5448 2567 5500 2576
rect 5448 2533 5475 2567
rect 5475 2533 5500 2567
rect 5448 2524 5500 2533
rect 5632 2567 5684 2576
rect 5632 2533 5641 2567
rect 5641 2533 5675 2567
rect 5675 2533 5684 2567
rect 5632 2524 5684 2533
rect 6552 2592 6604 2644
rect 7840 2592 7892 2644
rect 8576 2592 8628 2644
rect 8024 2524 8076 2576
rect 8116 2567 8168 2576
rect 8116 2533 8125 2567
rect 8125 2533 8159 2567
rect 8159 2533 8168 2567
rect 8116 2524 8168 2533
rect 8668 2524 8720 2576
rect 6184 2388 6236 2440
rect 7380 2456 7432 2508
rect 8208 2456 8260 2508
rect 6644 2388 6696 2440
rect 8484 2388 8536 2440
rect 7472 2320 7524 2372
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 5264 2295 5316 2304
rect 5264 2261 5273 2295
rect 5273 2261 5307 2295
rect 5307 2261 5316 2295
rect 5264 2252 5316 2261
rect 5908 2252 5960 2304
rect 6000 2295 6052 2304
rect 6000 2261 6009 2295
rect 6009 2261 6043 2295
rect 6043 2261 6052 2295
rect 6000 2252 6052 2261
rect 6460 2252 6512 2304
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 7748 2252 7800 2304
rect 8392 2252 8444 2304
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 4804 2048 4856 2100
rect 6000 2048 6052 2100
rect 6552 2048 6604 2100
rect 7748 2091 7800 2100
rect 7748 2057 7757 2091
rect 7757 2057 7791 2091
rect 7791 2057 7800 2091
rect 7748 2048 7800 2057
rect 8208 2048 8260 2100
rect 4252 1912 4304 1964
rect 4896 1887 4948 1896
rect 4896 1853 4905 1887
rect 4905 1853 4939 1887
rect 4939 1853 4948 1887
rect 4896 1844 4948 1853
rect 5264 1887 5316 1896
rect 5264 1853 5298 1887
rect 5298 1853 5316 1887
rect 5264 1844 5316 1853
rect 6460 1887 6512 1896
rect 6460 1853 6469 1887
rect 6469 1853 6503 1887
rect 6503 1853 6512 1887
rect 6460 1844 6512 1853
rect 6644 1887 6696 1896
rect 6644 1853 6653 1887
rect 6653 1853 6687 1887
rect 6687 1853 6696 1887
rect 6644 1844 6696 1853
rect 9772 1887 9824 1896
rect 9772 1853 9781 1887
rect 9781 1853 9815 1887
rect 9815 1853 9824 1887
rect 9772 1844 9824 1853
rect 3516 1776 3568 1828
rect 6184 1776 6236 1828
rect 7104 1819 7156 1828
rect 7104 1785 7131 1819
rect 7131 1785 7156 1819
rect 7104 1776 7156 1785
rect 7288 1819 7340 1828
rect 7288 1785 7297 1819
rect 7297 1785 7331 1819
rect 7331 1785 7340 1819
rect 7288 1776 7340 1785
rect 7840 1776 7892 1828
rect 4160 1708 4212 1760
rect 6920 1751 6972 1760
rect 6920 1717 6929 1751
rect 6929 1717 6963 1751
rect 6963 1717 6972 1751
rect 6920 1708 6972 1717
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 5908 1504 5960 1556
rect 6644 1504 6696 1556
rect 4160 1436 4212 1488
rect 4896 1436 4948 1488
rect 4252 1411 4304 1420
rect 4252 1377 4261 1411
rect 4261 1377 4295 1411
rect 4295 1377 4304 1411
rect 4252 1368 4304 1377
rect 6000 1411 6052 1420
rect 6000 1377 6009 1411
rect 6009 1377 6043 1411
rect 6043 1377 6052 1411
rect 6000 1368 6052 1377
rect 6184 1411 6236 1420
rect 5448 1300 5500 1352
rect 6184 1377 6193 1411
rect 6193 1377 6227 1411
rect 6227 1377 6236 1411
rect 6184 1368 6236 1377
rect 6920 1436 6972 1488
rect 6460 1368 6512 1420
rect 9772 1300 9824 1352
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 2688 892 2740 944
rect 8116 892 8168 944
rect 2964 799 3016 808
rect 2964 765 2973 799
rect 2973 765 3007 799
rect 3007 765 3016 799
rect 2964 756 3016 765
rect 7656 756 7708 808
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
<< metal2 >>
rect 386 10050 442 10850
rect 1214 10050 1270 10850
rect 2042 10050 2098 10850
rect 2870 10050 2926 10850
rect 3698 10050 3754 10850
rect 4526 10050 4582 10850
rect 5354 10050 5410 10850
rect 6182 10050 6238 10850
rect 7010 10050 7066 10850
rect 7838 10050 7894 10850
rect 8666 10050 8722 10850
rect 9494 10050 9550 10850
rect 10322 10050 10378 10850
rect 400 8430 428 10050
rect 1228 9602 1256 10050
rect 1044 9574 1256 9602
rect 1044 9042 1072 9574
rect 1124 9444 1176 9450
rect 1124 9386 1176 9392
rect 1216 9444 1268 9450
rect 1216 9386 1268 9392
rect 1032 9036 1084 9042
rect 1032 8978 1084 8984
rect 1136 8634 1164 9386
rect 1228 8974 1256 9386
rect 1216 8968 1268 8974
rect 1216 8910 1268 8916
rect 1124 8628 1176 8634
rect 1124 8570 1176 8576
rect 1228 8498 1256 8910
rect 1216 8492 1268 8498
rect 1216 8434 1268 8440
rect 388 8424 440 8430
rect 388 8366 440 8372
rect 1228 7954 1256 8434
rect 2056 8362 2084 10050
rect 2884 9602 2912 10050
rect 3712 10010 3740 10050
rect 3528 9982 3740 10010
rect 2884 9574 3004 9602
rect 2976 9518 3004 9574
rect 3528 9518 3556 9982
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 4540 9722 4568 10050
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 2332 8022 2360 9318
rect 3252 9110 3280 9318
rect 3240 9104 3292 9110
rect 3240 9046 3292 9052
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 2700 7954 2728 8774
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 1216 7948 1268 7954
rect 1216 7890 1268 7896
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 1228 6866 1256 7890
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2792 7410 2820 7686
rect 3068 7410 3096 8230
rect 3528 8022 3556 9318
rect 4172 8974 4200 9454
rect 4322 9276 4630 9285
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 4172 8294 4200 8910
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 3516 8016 3568 8022
rect 3516 7958 3568 7964
rect 4172 7954 4200 8230
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 2044 7336 2096 7342
rect 2044 7278 2096 7284
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 1308 7200 1360 7206
rect 1308 7142 1360 7148
rect 1216 6860 1268 6866
rect 1216 6802 1268 6808
rect 940 6248 992 6254
rect 940 6190 992 6196
rect 952 4622 980 6190
rect 1320 6186 1348 7142
rect 1308 6180 1360 6186
rect 1308 6122 1360 6128
rect 2056 5914 2084 7278
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2424 5914 2452 7142
rect 2516 6798 2544 7278
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2516 6322 2544 6734
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2240 5302 2268 5646
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1504 4758 1532 4966
rect 1492 4752 1544 4758
rect 1492 4694 1544 4700
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 1308 4480 1360 4486
rect 1308 4422 1360 4428
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 1320 4078 1348 4422
rect 2332 4214 2360 4422
rect 2320 4208 2372 4214
rect 2320 4150 2372 4156
rect 2792 4146 2820 4558
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 1308 4072 1360 4078
rect 1308 4014 1360 4020
rect 1320 3670 1348 4014
rect 1308 3664 1360 3670
rect 1308 3606 1360 3612
rect 2688 944 2740 950
rect 2688 886 2740 892
rect 2700 800 2728 886
rect 2976 814 3004 6598
rect 3068 5914 3096 6598
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3252 5574 3280 6190
rect 3344 5846 3372 7686
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 4172 7324 4200 7890
rect 4264 7478 4292 8774
rect 5368 8430 5396 10050
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5644 9178 5672 9454
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5736 8634 5764 8978
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 5092 8090 5120 8366
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4252 7336 4304 7342
rect 4172 7296 4252 7324
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6458 3464 6802
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3528 6254 3556 7142
rect 4172 6866 4200 7296
rect 4252 7278 4304 7284
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 4816 6934 4844 7142
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 5000 6866 5028 7686
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4264 5914 4292 6190
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3068 2922 3096 4422
rect 3160 4282 3188 5034
rect 3252 4486 3280 5510
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 4264 5302 4292 5850
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 4252 5296 4304 5302
rect 4252 5238 4304 5244
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3160 4078 3188 4218
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3252 3670 3280 4422
rect 3436 4162 3464 5238
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4540 5114 4568 5714
rect 4724 5710 4752 6258
rect 5552 5846 5580 8298
rect 5644 7954 5672 8502
rect 5828 8498 5856 9318
rect 6196 8498 6224 10050
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5736 7342 5764 8230
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 6472 6866 6500 8230
rect 6564 7954 6592 9318
rect 6840 9110 6868 9454
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6748 8634 6776 8978
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6840 7954 6868 9046
rect 7024 9042 7052 10050
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7300 8498 7328 8774
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6840 7410 6868 7890
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6840 6934 6868 7346
rect 7116 7342 7144 8230
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3528 4282 3556 4966
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3436 4134 3556 4162
rect 4172 4146 4200 4626
rect 4264 4214 4292 5102
rect 4540 5098 4752 5114
rect 4528 5092 4752 5098
rect 4580 5086 4752 5092
rect 4528 5034 4580 5040
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3160 3194 3188 3538
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3436 2938 3464 4134
rect 3528 4078 3556 4134
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4448 4078 4476 4626
rect 4724 4570 4752 5086
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 4690 5396 4966
rect 5552 4758 5580 5782
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 5736 5166 5764 5578
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5828 4865 5856 5170
rect 6104 5166 6132 6598
rect 7024 6322 7052 7142
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6748 5302 6776 5510
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6748 5166 6776 5238
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 5814 4856 5870 4865
rect 5814 4791 5870 4800
rect 5540 4752 5592 4758
rect 5446 4720 5502 4729
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 5356 4684 5408 4690
rect 5540 4694 5592 4700
rect 5446 4655 5448 4664
rect 5356 4626 5408 4632
rect 5500 4655 5502 4664
rect 5448 4626 5500 4632
rect 4632 4542 4752 4570
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4632 3942 4660 4542
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 3528 3194 3556 3878
rect 4172 3738 4200 3878
rect 4322 3836 4630 3845
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 4172 3210 4200 3538
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4080 3194 4200 3210
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 4068 3188 4200 3194
rect 4120 3182 4200 3188
rect 4068 3130 4120 3136
rect 3436 2922 3556 2938
rect 3056 2916 3108 2922
rect 3436 2916 3568 2922
rect 3436 2910 3516 2916
rect 3056 2858 3108 2864
rect 3516 2858 3568 2864
rect 3528 1834 3556 2858
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 4264 1970 4292 3334
rect 4724 2854 4752 4422
rect 4816 4282 4844 4626
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 5368 4146 5396 4626
rect 6104 4554 6132 5102
rect 6840 5098 6868 5306
rect 7024 5166 7052 6258
rect 7116 6254 7144 6598
rect 7300 6322 7328 7686
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7012 5160 7064 5166
rect 6932 5120 7012 5148
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4816 2990 4844 3878
rect 5092 3738 5120 4014
rect 5644 3942 5672 4422
rect 6288 4078 6316 4422
rect 6472 4214 6500 4966
rect 6564 4690 6592 4966
rect 6734 4856 6790 4865
rect 6734 4791 6790 4800
rect 6748 4758 6776 4791
rect 6736 4752 6788 4758
rect 6736 4694 6788 4700
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6564 4282 6592 4626
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 4816 2514 4844 2926
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 5644 2582 5672 2858
rect 6840 2774 6868 5034
rect 6932 4826 6960 5120
rect 7012 5102 7064 5108
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6918 4720 6974 4729
rect 7116 4672 7144 6054
rect 7300 5778 7328 6258
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 6974 4664 7144 4672
rect 6918 4655 6920 4664
rect 6972 4644 7144 4664
rect 6920 4626 6972 4632
rect 7208 4282 7236 5102
rect 7392 4690 7420 9318
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7668 7954 7696 8774
rect 7760 8634 7788 9386
rect 7852 9194 7880 10050
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 7852 9166 7972 9194
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7852 8362 7880 8978
rect 7944 8430 7972 9166
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 6866 8064 7686
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7944 6458 7972 6598
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7484 4826 7512 5782
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7300 4078 7328 4626
rect 7392 4146 7420 4626
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7300 3738 7328 4014
rect 7484 4010 7512 4626
rect 7576 4282 7604 4626
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 6564 2746 6868 2774
rect 6564 2650 6592 2746
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4816 2394 4844 2450
rect 4816 2366 4936 2394
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4816 2106 4844 2246
rect 4804 2100 4856 2106
rect 4804 2042 4856 2048
rect 4252 1964 4304 1970
rect 4252 1906 4304 1912
rect 3516 1828 3568 1834
rect 3516 1770 3568 1776
rect 4160 1760 4212 1766
rect 4160 1702 4212 1708
rect 4172 1494 4200 1702
rect 4160 1488 4212 1494
rect 4160 1430 4212 1436
rect 4264 1426 4292 1906
rect 4908 1902 4936 2366
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 5276 1902 5304 2246
rect 4896 1896 4948 1902
rect 4896 1838 4948 1844
rect 5264 1896 5316 1902
rect 5264 1838 5316 1844
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 4908 1494 4936 1838
rect 4896 1488 4948 1494
rect 4896 1430 4948 1436
rect 4252 1420 4304 1426
rect 4252 1362 4304 1368
rect 5460 1358 5488 2518
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 5920 1562 5948 2246
rect 6012 2106 6040 2246
rect 6000 2100 6052 2106
rect 6000 2042 6052 2048
rect 5908 1556 5960 1562
rect 5908 1498 5960 1504
rect 6012 1426 6040 2042
rect 6196 1834 6224 2382
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6472 1902 6500 2246
rect 6564 2106 6592 2586
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6552 2100 6604 2106
rect 6552 2042 6604 2048
rect 6656 1902 6684 2382
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 6460 1896 6512 1902
rect 6460 1838 6512 1844
rect 6644 1896 6696 1902
rect 6644 1838 6696 1844
rect 6184 1828 6236 1834
rect 6184 1770 6236 1776
rect 6196 1426 6224 1770
rect 6472 1426 6500 1838
rect 6656 1562 6684 1838
rect 7116 1834 7144 2246
rect 7300 1834 7328 2858
rect 7392 2514 7420 3538
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 7484 2378 7512 3946
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 7104 1828 7156 1834
rect 7104 1770 7156 1776
rect 7288 1828 7340 1834
rect 7288 1770 7340 1776
rect 6920 1760 6972 1766
rect 6920 1702 6972 1708
rect 6644 1556 6696 1562
rect 6644 1498 6696 1504
rect 6932 1494 6960 1702
rect 6920 1488 6972 1494
rect 6920 1430 6972 1436
rect 6000 1420 6052 1426
rect 6000 1362 6052 1368
rect 6184 1420 6236 1426
rect 6184 1362 6236 1368
rect 6460 1420 6512 1426
rect 6460 1362 6512 1368
rect 5448 1352 5500 1358
rect 5448 1294 5500 1300
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 7668 814 7696 6258
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7760 4826 7788 5102
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7852 4622 7880 5850
rect 7944 5778 7972 6394
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 8128 5642 8156 9318
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8404 7546 8432 7822
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8036 4690 8064 5510
rect 8220 5166 8248 7142
rect 8496 6866 8524 9386
rect 8680 9042 8708 10050
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9416 7274 9444 8774
rect 9508 7954 9536 10050
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9968 8974 9996 9454
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9968 8430 9996 8910
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9692 8090 9720 8298
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9508 6934 9536 7686
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8680 5778 8708 6598
rect 9784 6322 9812 7278
rect 9968 6866 9996 8366
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9508 5914 9536 6122
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8864 5234 8892 5646
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 8036 3602 8064 4422
rect 8220 3670 8248 4966
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 7760 3126 7788 3538
rect 7748 3120 7800 3126
rect 7748 3062 7800 3068
rect 7852 2650 7880 3538
rect 8036 3398 8064 3538
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 8220 3058 8248 3606
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8312 3194 8340 3538
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8116 2916 8168 2922
rect 8116 2858 8168 2864
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 2106 7788 2246
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 7852 1834 7880 2586
rect 8036 2582 8064 2790
rect 8128 2582 8156 2858
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 8220 2514 8248 2858
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8220 2106 8248 2450
rect 8404 2310 8432 3402
rect 8496 2446 8524 5170
rect 8864 4282 8892 5170
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8680 3602 8708 3674
rect 8956 3670 8984 5510
rect 9784 4758 9812 6258
rect 10336 5846 10364 10050
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9876 5370 9904 5714
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 9048 3738 9076 3946
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 9232 3602 9260 4218
rect 9784 4078 9812 4694
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8588 2650 8616 2858
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8680 2582 8708 3538
rect 9140 3194 9168 3538
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9784 2990 9812 4014
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 9784 1902 9812 2926
rect 9772 1896 9824 1902
rect 9772 1838 9824 1844
rect 7840 1828 7892 1834
rect 7840 1770 7892 1776
rect 9784 1358 9812 1838
rect 9772 1352 9824 1358
rect 9772 1294 9824 1300
rect 8116 944 8168 950
rect 8116 886 8168 892
rect 2964 808 3016 814
rect 2686 0 2742 800
rect 2964 750 3016 756
rect 7656 808 7708 814
rect 8128 800 8156 886
rect 7656 750 7708 756
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
rect 8114 0 8170 800
<< via2 >>
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 5814 4800 5870 4856
rect 5446 4684 5502 4720
rect 5446 4664 5448 4684
rect 5448 4664 5500 4684
rect 5500 4664 5502 4684
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 6734 4800 6790 4856
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 6918 4684 6974 4720
rect 6918 4664 6920 4684
rect 6920 4664 6972 4684
rect 6972 4664 6974 4684
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
<< metal3 >>
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 5809 4858 5875 4861
rect 6729 4858 6795 4861
rect 5809 4856 6795 4858
rect 5809 4800 5814 4856
rect 5870 4800 6734 4856
rect 6790 4800 6795 4856
rect 5809 4798 6795 4800
rect 5809 4795 5875 4798
rect 6729 4795 6795 4798
rect 5441 4722 5507 4725
rect 6913 4722 6979 4725
rect 5441 4720 6979 4722
rect 5441 4664 5446 4720
rect 5502 4664 6918 4720
rect 6974 4664 6979 4720
rect 5441 4662 6979 4664
rect 5441 4659 5507 4662
rect 6913 4659 6979 4662
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 4318 3775 4634 3776
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
<< via3 >>
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
<< metal4 >>
rect 3656 9824 3976 9840
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 9280 4636 9840
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4316 8192 4636 9216
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
use sky130_fd_sc_hd__inv_2  _053_
timestamp 28801
transform 1 0 5152 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _054_
timestamp 28801
transform -1 0 5152 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _055_
timestamp 28801
transform 1 0 7912 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp 28801
transform 1 0 7636 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 28801
transform -1 0 7452 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 28801
transform -1 0 8372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059_
timestamp 28801
transform -1 0 9936 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _060_
timestamp 28801
transform 1 0 3496 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _061_
timestamp 28801
transform 1 0 2668 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _062_
timestamp 28801
transform 1 0 6072 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__xor2_1  _063_
timestamp 28801
transform -1 0 9016 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _064_
timestamp 28801
transform 1 0 4324 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _065_
timestamp 28801
transform 1 0 4048 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _066_
timestamp 28801
transform 1 0 7084 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _067_
timestamp 28801
transform 1 0 6532 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _068_
timestamp 28801
transform 1 0 5704 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _069_
timestamp 28801
transform -1 0 8924 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _070_
timestamp 28801
transform -1 0 7084 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _071_
timestamp 28801
transform 1 0 6992 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _072_
timestamp 28801
transform -1 0 5704 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _073_
timestamp 28801
transform 1 0 6348 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _074_
timestamp 28801
transform 1 0 7268 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _075_
timestamp 28801
transform -1 0 2852 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _076_
timestamp 28801
transform 1 0 1656 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _077_
timestamp 28801
transform -1 0 2024 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _078_
timestamp 28801
transform 1 0 3220 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _079_
timestamp 28801
transform -1 0 3128 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _080_
timestamp 28801
transform -1 0 3680 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _081_
timestamp 28801
transform 1 0 3680 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _082_
timestamp 28801
transform 1 0 2484 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _083_
timestamp 28801
transform -1 0 3680 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _084_
timestamp 28801
transform 1 0 4232 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _085_
timestamp 28801
transform -1 0 4692 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _086_
timestamp 28801
transform 1 0 4600 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _087_
timestamp 28801
transform -1 0 4416 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _088_
timestamp 28801
transform -1 0 4968 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _089_
timestamp 28801
transform -1 0 4968 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _090_
timestamp 28801
transform 1 0 4048 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _091_
timestamp 28801
transform 1 0 5796 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 28801
transform 1 0 6348 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _093_
timestamp 28801
transform 1 0 5796 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _094_
timestamp 28801
transform -1 0 5704 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _095_
timestamp 28801
transform 1 0 6440 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _096_
timestamp 28801
transform 1 0 6256 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _097_
timestamp 28801
transform -1 0 7268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _098_
timestamp 28801
transform -1 0 7360 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _099_
timestamp 28801
transform -1 0 8004 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _100_
timestamp 28801
transform 1 0 7268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _101_
timestamp 28801
transform 1 0 7544 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _102_
timestamp 28801
transform 1 0 7820 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _103_
timestamp 28801
transform -1 0 8280 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 28801
transform -1 0 7820 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _105_
timestamp 28801
transform 1 0 8096 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _106_
timestamp 28801
transform 1 0 9108 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _107_
timestamp 28801
transform -1 0 9108 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _108_
timestamp 28801
transform 1 0 920 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _109_
timestamp 28801
transform 1 0 920 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _110_
timestamp 28801
transform 1 0 1288 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _111_
timestamp 28801
transform 1 0 2392 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _112_
timestamp 28801
transform 1 0 3864 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _113_
timestamp 28801
transform 1 0 4232 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _114_
timestamp 28801
transform 1 0 4968 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _115_
timestamp 28801
transform -1 0 8280 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _116_
timestamp 28801
transform -1 0 9844 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _117_
timestamp 28801
transform -1 0 9936 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _118_
timestamp 28801
transform -1 0 9936 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _119_
timestamp 28801
transform 1 0 828 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _120_
timestamp 28801
transform 1 0 1104 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _121_
timestamp 28801
transform -1 0 10028 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _122_
timestamp 28801
transform 1 0 1196 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _123_
timestamp 28801
transform 1 0 1288 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _124_
timestamp 28801
transform 1 0 1656 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _125_
timestamp 28801
transform 1 0 2760 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _126_
timestamp 28801
transform 1 0 3404 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _127_
timestamp 28801
transform 1 0 4140 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _128_
timestamp 28801
transform 1 0 4232 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _129_
timestamp 28801
transform 1 0 5888 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _130_
timestamp 28801
transform 1 0 7360 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _131_
timestamp 28801
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _132_
timestamp 28801
transform -1 0 9844 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _133_
timestamp 28801
transform 1 0 2852 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _134_
timestamp 28801
transform 1 0 3220 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _135_
timestamp 28801
transform 1 0 4140 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _136_
timestamp 28801
transform 1 0 4876 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _137_
timestamp 28801
transform 1 0 5796 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _138_
timestamp 28801
transform 1 0 5796 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _139_
timestamp 28801
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _140_
timestamp 28801
transform 1 0 8372 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _141_
timestamp 28801
transform -1 0 9844 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _142_
timestamp 28801
transform -1 0 10028 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK
timestamp 28801
transform -1 0 7636 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_CLK
timestamp 28801
transform -1 0 4600 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_CLK
timestamp 28801
transform 1 0 3220 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_CLK
timestamp 28801
transform 1 0 8188 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_CLK
timestamp 28801
transform 1 0 7820 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp 28801
transform -1 0 7820 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636997256
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_15
timestamp 28801
transform 1 0 1932 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_23
timestamp 28801
transform 1 0 2668 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 28801
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636997256
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636997256
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 28801
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636997256
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636997256
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 28801
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_89
timestamp 1636997256
transform 1 0 8740 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_101
timestamp 28801
transform 1 0 9844 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636997256
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636997256
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636997256
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_39
timestamp 28801
transform 1 0 4140 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_66
timestamp 28801
transform 1 0 6624 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_84
timestamp 1636997256
transform 1 0 8280 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_96
timestamp 28801
transform 1 0 9384 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_102
timestamp 28801
transform 1 0 9936 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636997256
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636997256
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 28801
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 28801
transform 1 0 3220 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_37
timestamp 28801
transform 1 0 3956 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_74
timestamp 28801
transform 1 0 7360 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 28801
transform 1 0 8004 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_101
timestamp 28801
transform 1 0 9844 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636997256
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636997256
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636997256
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_39
timestamp 28801
transform 1 0 4140 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_48
timestamp 28801
transform 1 0 4968 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_69
timestamp 28801
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_81
timestamp 28801
transform 1 0 8004 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_87
timestamp 1636997256
transform 1 0 8556 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_99
timestamp 28801
transform 1 0 9660 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636997256
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636997256
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 28801
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_34
timestamp 28801
transform 1 0 3680 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_45
timestamp 1636997256
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_57
timestamp 1636997256
transform 1 0 5796 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_69
timestamp 28801
transform 1 0 6900 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 28801
transform 1 0 8372 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_102
timestamp 28801
transform 1 0 9936 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636997256
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_15
timestamp 28801
transform 1 0 1932 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_19
timestamp 28801
transform 1 0 2300 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 28801
transform 1 0 5336 0 -1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636997256
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_69
timestamp 28801
transform 1 0 6900 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_75
timestamp 28801
transform 1 0 7452 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_98
timestamp 28801
transform 1 0 9568 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_102
timestamp 28801
transform 1 0 9936 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 28801
transform 1 0 828 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_7
timestamp 28801
transform 1 0 1196 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_24
timestamp 28801
transform 1 0 2760 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_39
timestamp 28801
transform 1 0 4140 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_53
timestamp 28801
transform 1 0 5428 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_61
timestamp 28801
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 28801
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 28801
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 28801
transform 1 0 8372 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_102
timestamp 28801
transform 1 0 9936 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 28801
transform 1 0 828 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_20
timestamp 28801
transform 1 0 2392 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_47
timestamp 28801
transform 1 0 4876 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 28801
transform 1 0 5796 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_61
timestamp 28801
transform 1 0 6164 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_79
timestamp 28801
transform 1 0 7820 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_3
timestamp 28801
transform 1 0 828 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_9
timestamp 28801
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_16
timestamp 28801
transform 1 0 2024 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_25
timestamp 28801
transform 1 0 2852 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_34
timestamp 28801
transform 1 0 3680 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_45
timestamp 28801
transform 1 0 4692 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_53
timestamp 28801
transform 1 0 5428 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_80
timestamp 28801
transform 1 0 7912 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_92
timestamp 28801
transform 1 0 9016 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 28801
transform 1 0 828 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_11
timestamp 28801
transform 1 0 1564 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_21
timestamp 28801
transform 1 0 2484 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_48
timestamp 28801
transform 1 0 4968 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_83
timestamp 28801
transform 1 0 8188 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_102
timestamp 28801
transform 1 0 9936 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 28801
transform 1 0 828 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_45
timestamp 1636997256
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_57
timestamp 28801
transform 1 0 5796 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 28801
transform 1 0 8004 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_101
timestamp 28801
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_3
timestamp 28801
transform 1 0 828 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_35
timestamp 28801
transform 1 0 3772 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 28801
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_73
timestamp 28801
transform 1 0 7268 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 28801
transform 1 0 828 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_9
timestamp 28801
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_18
timestamp 28801
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25
timestamp 28801
transform 1 0 2852 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 28801
transform 1 0 3220 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_38
timestamp 28801
transform 1 0 4048 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_63
timestamp 28801
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_67
timestamp 28801
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_101
timestamp 28801
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_3
timestamp 28801
transform 1 0 828 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_22
timestamp 28801
transform 1 0 2576 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_47
timestamp 28801
transform 1 0 4876 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_73
timestamp 28801
transform 1 0 7268 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_101
timestamp 28801
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_6
timestamp 28801
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_71
timestamp 28801
transform 1 0 7084 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 28801
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 28801
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 28801
transform 1 0 828 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 28801
transform 1 0 5796 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_77
timestamp 28801
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_102
timestamp 28801
transform 1 0 9936 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 28801
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_32
timestamp 28801
transform 1 0 3496 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_55
timestamp 28801
transform 1 0 5612 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_57
timestamp 28801
transform 1 0 5796 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_66
timestamp 28801
transform 1 0 6624 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_101
timestamp 28801
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 28801
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 28801
transform 1 0 5060 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 28801
transform -1 0 7912 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 28801
transform 1 0 7820 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 28801
transform -1 0 3036 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 28801
transform 1 0 4140 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 28801
transform 1 0 5888 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 28801
transform 1 0 3312 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 28801
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 28801
transform 1 0 2668 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 28801
transform -1 0 5704 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 28801
transform 1 0 8924 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 28801
transform 1 0 2392 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 28801
transform -1 0 2208 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 28801
transform 1 0 9292 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 28801
transform -1 0 2852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 28801
transform -1 0 9844 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 28801
transform -1 0 1288 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 28801
transform -1 0 1656 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 28801
transform 1 0 3220 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 28801
transform 1 0 3588 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 28801
transform -1 0 4140 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 28801
transform 1 0 6532 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 28801
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 28801
transform -1 0 7636 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 28801
transform 1 0 7912 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 28801
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 28801
transform -1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output13
timestamp 28801
transform 1 0 2760 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 28801
transform 1 0 8372 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_17
timestamp 28801
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 28801
transform -1 0 10304 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_18
timestamp 28801
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 28801
transform -1 0 10304 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_19
timestamp 28801
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 28801
transform -1 0 10304 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_20
timestamp 28801
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 28801
transform -1 0 10304 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_21
timestamp 28801
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 28801
transform -1 0 10304 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_22
timestamp 28801
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 28801
transform -1 0 10304 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_23
timestamp 28801
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 28801
transform -1 0 10304 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_24
timestamp 28801
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 28801
transform -1 0 10304 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_25
timestamp 28801
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 28801
transform -1 0 10304 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_26
timestamp 28801
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 28801
transform -1 0 10304 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_27
timestamp 28801
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 28801
transform -1 0 10304 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_28
timestamp 28801
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 28801
transform -1 0 10304 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_29
timestamp 28801
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 28801
transform -1 0 10304 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_30
timestamp 28801
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 28801
transform -1 0 10304 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_31
timestamp 28801
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 28801
transform -1 0 10304 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_32
timestamp 28801
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 28801
transform -1 0 10304 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_33
timestamp 28801
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 28801
transform -1 0 10304 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp 28801
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp 28801
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp 28801
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_37
timestamp 28801
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_38
timestamp 28801
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_39
timestamp 28801
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_40
timestamp 28801
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_41
timestamp 28801
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_42
timestamp 28801
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_43
timestamp 28801
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_44
timestamp 28801
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_45
timestamp 28801
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_46
timestamp 28801
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_47
timestamp 28801
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_48
timestamp 28801
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_49
timestamp 28801
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_50
timestamp 28801
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_51
timestamp 28801
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_52
timestamp 28801
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_53
timestamp 28801
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_54
timestamp 28801
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_55
timestamp 28801
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_56
timestamp 28801
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_57
timestamp 28801
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_58
timestamp 28801
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_59
timestamp 28801
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_60
timestamp 28801
transform 1 0 5704 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_61
timestamp 28801
transform 1 0 8280 0 1 9248
box -38 -48 130 592
<< labels >>
flabel metal2 s 10322 10050 10378 10850 0 FreeSans 224 90 0 0 CLK
port 0 nsew signal input
flabel metal2 s 2686 0 2742 800 0 FreeSans 224 90 0 0 CLK_OUT
port 1 nsew signal output
flabel metal2 s 9494 10050 9550 10850 0 FreeSans 224 90 0 0 ENABLE
port 2 nsew signal input
flabel metal2 s 1214 10050 1270 10850 0 FreeSans 224 90 0 0 N[0]
port 3 nsew signal input
flabel metal2 s 2042 10050 2098 10850 0 FreeSans 224 90 0 0 N[1]
port 4 nsew signal input
flabel metal2 s 2870 10050 2926 10850 0 FreeSans 224 90 0 0 N[2]
port 5 nsew signal input
flabel metal2 s 3698 10050 3754 10850 0 FreeSans 224 90 0 0 N[3]
port 6 nsew signal input
flabel metal2 s 4526 10050 4582 10850 0 FreeSans 224 90 0 0 N[4]
port 7 nsew signal input
flabel metal2 s 5354 10050 5410 10850 0 FreeSans 224 90 0 0 N[5]
port 8 nsew signal input
flabel metal2 s 6182 10050 6238 10850 0 FreeSans 224 90 0 0 N[6]
port 9 nsew signal input
flabel metal2 s 7010 10050 7066 10850 0 FreeSans 224 90 0 0 N[7]
port 10 nsew signal input
flabel metal2 s 7838 10050 7894 10850 0 FreeSans 224 90 0 0 N[8]
port 11 nsew signal input
flabel metal2 s 8666 10050 8722 10850 0 FreeSans 224 90 0 0 N[9]
port 12 nsew signal input
flabel metal2 s 386 10050 442 10850 0 FreeSans 224 90 0 0 RESETn
port 13 nsew signal input
flabel metal4 s 4316 496 4636 9840 0 FreeSans 1920 90 0 0 VGND
port 14 nsew ground bidirectional
flabel metal4 s 3656 496 3976 9840 0 FreeSans 1920 90 0 0 VPWR
port 15 nsew power bidirectional
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 temp
port 16 nsew signal output
rlabel metal1 5428 9248 5428 9248 0 VGND
rlabel metal1 5428 9792 5428 9792 0 VPWR
rlabel metal1 8970 5814 8970 5814 0 CLK
rlabel metal2 2714 840 2714 840 0 CLK_OUT
rlabel metal1 9568 7922 9568 7922 0 ENABLE
rlabel metal2 1058 9299 1058 9299 0 N[0]
rlabel metal1 1748 8398 1748 8398 0 N[1]
rlabel metal1 3220 9486 3220 9486 0 N[2]
rlabel metal1 3680 9486 3680 9486 0 N[3]
rlabel metal1 3910 9588 3910 9588 0 N[4]
rlabel metal1 6072 8398 6072 8398 0 N[5]
rlabel metal1 7038 8432 7038 8432 0 N[6]
rlabel metal1 7222 9010 7222 9010 0 N[7]
rlabel metal1 8050 8398 8050 8398 0 N[8]
rlabel metal1 9292 9010 9292 9010 0 N[9]
rlabel metal1 644 8398 644 8398 0 RESETn
rlabel metal1 1886 5882 1886 5882 0 _000_
rlabel metal1 1375 4726 1375 4726 0 _001_
rlabel metal1 3266 3944 3266 3944 0 _002_
rlabel metal1 3220 3162 3220 3162 0 _003_
rlabel metal1 4048 3162 4048 3162 0 _004_
rlabel metal1 4360 1462 4360 1462 0 _005_
rlabel via1 5285 1870 5285 1870 0 _006_
rlabel metal1 7456 1462 7456 1462 0 _007_
rlabel metal1 8744 1802 8744 1802 0 _008_
rlabel metal1 8556 2618 8556 2618 0 _009_
rlabel metal2 9062 3842 9062 3842 0 _010_
rlabel metal1 3910 4080 3910 4080 0 _011_
rlabel metal1 6532 4658 6532 4658 0 _012_
rlabel metal1 7843 4658 7843 4658 0 _013_
rlabel via1 6744 5134 6744 5134 0 _014_
rlabel metal2 7314 4352 7314 4352 0 _015_
rlabel metal1 6210 4590 6210 4590 0 _016_
rlabel viali 8819 3570 8819 3570 0 _017_
rlabel metal1 2415 5746 2415 5746 0 _018_
rlabel metal1 6578 5168 6578 5168 0 _019_
rlabel metal2 5750 5372 5750 5372 0 _020_
rlabel metal1 7130 4692 7130 4692 0 _021_
rlabel metal2 7774 4964 7774 4964 0 _022_
rlabel metal1 7314 5338 7314 5338 0 _023_
rlabel metal1 6440 4182 6440 4182 0 _024_
rlabel metal1 7038 4624 7038 4624 0 _025_
rlabel metal1 6440 4046 6440 4046 0 _026_
rlabel metal1 6854 3978 6854 3978 0 _027_
rlabel metal1 6210 3910 6210 3910 0 _028_
rlabel metal1 7084 4250 7084 4250 0 _029_
rlabel metal1 8418 3604 8418 3604 0 _030_
rlabel metal1 2300 5882 2300 5882 0 _031_
rlabel metal1 3496 4250 3496 4250 0 _032_
rlabel metal1 2530 4624 2530 4624 0 _033_
rlabel metal1 3818 3910 3818 3910 0 _034_
rlabel metal2 3082 3672 3082 3672 0 _035_
rlabel metal1 4876 2482 4876 2482 0 _036_
rlabel metal1 4370 3162 4370 3162 0 _037_
rlabel metal1 4454 2822 4454 2822 0 _038_
rlabel metal1 4554 2074 4554 2074 0 _039_
rlabel metal1 4432 1802 4432 1802 0 _040_
rlabel metal2 6486 2074 6486 2074 0 _041_
rlabel metal1 6210 1530 6210 1530 0 _042_
rlabel metal1 5658 1326 5658 1326 0 _043_
rlabel metal1 6992 2074 6992 2074 0 _044_
rlabel metal1 8004 2550 8004 2550 0 _045_
rlabel via1 7122 1802 7122 1802 0 _046_
rlabel metal2 7774 2176 7774 2176 0 _047_
rlabel metal1 7682 2618 7682 2618 0 _048_
rlabel metal1 8372 2278 8372 2278 0 _049_
rlabel metal1 8234 3094 8234 3094 0 _050_
rlabel metal1 8526 2550 8526 2550 0 _051_
rlabel metal1 8602 3502 8602 3502 0 _052_
rlabel metal2 4278 6052 4278 6052 0 a\[0\]
rlabel metal1 4646 6324 4646 6324 0 a\[1\]
rlabel metal2 6118 4828 6118 4828 0 a\[2\]
rlabel metal2 7038 6732 7038 6732 0 a\[3\]
rlabel metal1 5060 4726 5060 4726 0 clknet_0_CLK
rlabel metal1 2438 3604 2438 3604 0 clknet_2_0__leaf_CLK
rlabel metal1 1196 7922 1196 7922 0 clknet_2_1__leaf_CLK
rlabel metal2 9798 1598 9798 1598 0 clknet_2_2__leaf_CLK
rlabel metal2 9982 7616 9982 7616 0 clknet_2_3__leaf_CLK
rlabel metal1 2714 4114 2714 4114 0 counter\[0\]
rlabel metal1 4554 3910 4554 3910 0 counter\[1\]
rlabel metal1 4462 3978 4462 3978 0 counter\[2\]
rlabel metal2 5106 3876 5106 3876 0 counter\[3\]
rlabel metal1 6900 2346 6900 2346 0 counter\[4\]
rlabel metal1 6532 2618 6532 2618 0 counter\[5\]
rlabel metal1 6578 2448 6578 2448 0 counter\[6\]
rlabel metal1 8004 2482 8004 2482 0 counter\[7\]
rlabel metal1 8280 3162 8280 3162 0 counter\[8\]
rlabel metal1 9108 5202 9108 5202 0 counter\[9\]
rlabel metal1 3266 6732 3266 6732 0 enable
rlabel metal2 5658 8228 5658 8228 0 enable0
rlabel metal2 2714 8364 2714 8364 0 n0\[0\]
rlabel metal1 3220 7378 3220 7378 0 n0\[1\]
rlabel metal1 4186 7412 4186 7412 0 n0\[2\]
rlabel metal1 4968 8058 4968 8058 0 n0\[3\]
rlabel metal2 5842 8908 5842 8908 0 n0\[4\]
rlabel metal2 5658 9316 5658 9316 0 n0\[5\]
rlabel metal1 7544 8466 7544 8466 0 n0\[6\]
rlabel metal1 8004 6834 8004 6834 0 n0\[7\]
rlabel metal1 8970 5644 8970 5644 0 n0\[8\]
rlabel metal2 8418 7684 8418 7684 0 n0\[9\]
rlabel metal1 7590 6630 7590 6630 0 n\[4\]
rlabel metal2 7314 7004 7314 7004 0 n\[5\]
rlabel metal1 8510 5134 8510 5134 0 n\[6\]
rlabel metal2 7406 7004 7406 7004 0 n\[7\]
rlabel viali 6854 4659 6854 4659 0 n\[8\]
rlabel metal2 8694 6188 8694 6188 0 n\[9\]
rlabel metal1 9752 8058 9752 8058 0 net1
rlabel metal1 7866 8602 7866 8602 0 net10
rlabel metal1 9480 7242 9480 7242 0 net11
rlabel metal1 1104 8602 1104 8602 0 net12
rlabel metal1 2852 6630 2852 6630 0 net13
rlabel metal1 8050 782 8050 782 0 net14
rlabel metal2 2254 5474 2254 5474 0 net15
rlabel metal1 9618 6902 9618 6902 0 net16
rlabel metal1 5469 7310 5469 7310 0 net17
rlabel via1 7125 7310 7125 7310 0 net18
rlabel metal2 8510 8126 8510 8126 0 net19
rlabel metal1 1416 9010 1416 9010 0 net2
rlabel metal1 1881 7990 1881 7990 0 net20
rlabel metal1 4641 6902 4641 6902 0 net21
rlabel metal1 6343 7922 6343 7922 0 net22
rlabel via1 3537 6222 3537 6222 0 net23
rlabel metal1 6297 6834 6297 6834 0 net24
rlabel metal1 3261 5814 3261 5814 0 net25
rlabel metal1 3358 6800 3358 6800 0 net26
rlabel metal1 9568 5882 9568 5882 0 net27
rlabel metal1 3266 6426 3266 6426 0 net28
rlabel metal1 1283 6154 1283 6154 0 net29
rlabel metal1 1778 8330 1778 8330 0 net3
rlabel metal1 9936 5338 9936 5338 0 net30
rlabel metal1 2070 5066 2070 5066 0 net31
rlabel metal1 3169 9078 3169 9078 0 net4
rlabel metal1 3618 7990 3618 7990 0 net5
rlabel metal1 4262 9418 4262 9418 0 net6
rlabel metal1 6164 8602 6164 8602 0 net7
rlabel metal1 6808 8602 6808 8602 0 net8
rlabel via1 7677 7922 7677 7922 0 net9
rlabel metal2 2530 6528 2530 6528 0 out
rlabel metal2 2806 7548 2806 7548 0 resetn
rlabel metal1 2507 9622 2507 9622 0 resetn0
rlabel metal2 8142 840 8142 840 0 temp
<< properties >>
string FIXED_BBOX 0 0 10866 10850
<< end >>
