magic
tech sky130A
magscale 1 2
timestamp 1717082902
<< metal1 >>
rect 26470 5040 26480 5430
rect 28820 5040 28830 5430
rect 26279 3650 26285 3760
rect 26395 3650 26401 3760
rect 28690 3076 31431 3186
rect 31321 2813 31431 3076
rect 26470 2690 26480 2800
rect 28810 2690 28820 2800
rect 31321 2697 31431 2703
<< via1 >>
rect 26480 5040 28820 5430
rect 26285 3650 26395 3760
rect 26480 2690 28810 2800
rect 31321 2703 31431 2813
<< metal2 >>
rect 26480 5430 28820 5440
rect 26480 5030 28820 5040
rect 26285 3760 26395 3766
rect 25736 3650 25745 3760
rect 25855 3650 26285 3760
rect 26285 3644 26395 3650
rect 26480 2800 28810 2810
rect 26480 2680 28810 2690
rect 31284 2675 31293 2842
rect 31460 2675 31469 2842
<< via2 >>
rect 26480 5040 28820 5430
rect 25745 3650 25855 3760
rect 26480 2690 28810 2800
rect 31293 2813 31460 2842
rect 31293 2703 31321 2813
rect 31321 2703 31431 2813
rect 31431 2703 31460 2813
rect 31293 2675 31460 2703
<< metal3 >>
rect 26470 5430 28830 5435
rect 190 5140 200 5430
rect 500 5140 26480 5430
rect 26470 5040 26480 5140
rect 28820 5040 28830 5430
rect 26470 5035 28830 5040
rect 25734 3645 25740 3765
rect 25850 3760 25860 3765
rect 25855 3650 25860 3760
rect 25850 3645 25860 3650
rect 9790 2660 9800 2950
rect 10100 2805 28810 2950
rect 10100 2800 28820 2805
rect 10100 2690 26480 2800
rect 28810 2690 28820 2800
rect 10100 2685 28820 2690
rect 10100 2660 28810 2685
rect 31269 2657 31275 2861
rect 31479 2657 31485 2861
<< via3 >>
rect 200 5140 500 5430
rect 25740 3760 25850 3765
rect 25740 3650 25745 3760
rect 25745 3650 25850 3760
rect 25740 3645 25850 3650
rect 9800 2660 10100 2950
rect 31275 2842 31479 2861
rect 31275 2675 31293 2842
rect 31293 2675 31460 2842
rect 31460 2675 31479 2842
rect 31275 2657 31479 2675
<< metal4 >>
rect 798 44460 858 45152
rect 1534 44800 1594 45152
rect 2270 44800 2330 45152
rect 3006 44800 3066 45152
rect 3742 44800 3802 45152
rect 4478 44800 4538 45152
rect 5214 44800 5274 45152
rect 5950 44800 6010 45152
rect 6686 44800 6746 45152
rect 7422 44800 7482 45152
rect 8158 44800 8218 45152
rect 8894 44800 8954 45152
rect 9630 44800 9690 45152
rect 10366 44800 10426 45152
rect 11102 44800 11162 45152
rect 11838 44800 11898 45152
rect 12574 44800 12634 45152
rect 13310 44800 13370 45152
rect 14046 44800 14106 45152
rect 14782 44800 14842 45152
rect 15518 44800 15578 45152
rect 16254 44800 16314 45152
rect 16990 44800 17050 45152
rect 1220 44460 17270 44800
rect 798 44400 17270 44460
rect 200 5431 500 44152
rect 1220 44110 17270 44400
rect 199 5430 501 5431
rect 199 5140 200 5430
rect 500 5140 501 5430
rect 199 5139 501 5140
rect 200 1000 500 5139
rect 9800 2951 10100 44110
rect 17726 3740 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 25739 3765 25851 3766
rect 25739 3740 25740 3765
rect 17726 3680 25740 3740
rect 25739 3645 25740 3680
rect 25850 3645 25851 3765
rect 25739 3644 25851 3645
rect 9799 2950 10101 2951
rect 9799 2660 9800 2950
rect 10100 2660 10101 2950
rect 9799 2659 10101 2660
rect 31274 2861 31480 2862
rect 9800 1000 10100 2659
rect 31274 2657 31275 2861
rect 31479 2657 31480 2861
rect 31274 2656 31480 2657
rect 31309 200 31446 2656
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 200
use ring_osc3  ring_osc3_0
timestamp 1717055118
transform -1 0 28010 0 1 3890
box -800 -1200 1730 1260
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
