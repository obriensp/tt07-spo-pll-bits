magic
tech sky130A
magscale 1 2
timestamp 1717029282
<< nwell >>
rect 1110 -1650 1620 -210
<< pwell >>
rect 1110 -2670 1620 -1660
<< metal1 >>
rect 1110 -320 1620 -210
rect 1150 -770 1300 -370
rect 1420 -770 1580 -320
rect 1150 -1030 1230 -770
rect 1260 -910 1460 -800
rect 1150 -1430 1300 -1030
rect 1420 -1430 1570 -1030
rect 1310 -1600 1410 -1470
rect 1110 -1710 1410 -1600
rect 1310 -1840 1410 -1710
rect 1470 -1600 1570 -1430
rect 1470 -1710 1620 -1600
rect 1470 -1870 1570 -1710
rect 1150 -2070 1300 -1870
rect 1420 -2070 1570 -1870
rect 1150 -2320 1230 -2070
rect 1260 -2290 1460 -2180
rect 1520 -2320 1580 -2270
rect 1150 -2520 1300 -2320
rect 1420 -2560 1580 -2320
rect 1110 -2670 1620 -2560
use sky130_fd_pr__nfet_01v8_46DABQ  sky130_fd_pr__nfet_01v8_46DABQ_0
timestamp 1717028433
transform 1 0 1361 0 1 -1941
box -241 -279 241 279
use sky130_fd_pr__nfet_01v8_TTGNW2  sky130_fd_pr__nfet_01v8_TTGNW2_0
timestamp 1717028433
transform 1 0 1361 0 1 -2391
box -241 -279 241 279
use sky130_fd_pr__pfet_01v8_5YCKZA  sky130_fd_pr__pfet_01v8_5YCKZA_0
timestamp 1717028433
transform 1 0 1361 0 1 -1266
box -241 -384 241 384
use sky130_fd_pr__pfet_01v8_38U2ME  sky130_fd_pr__pfet_01v8_38U2ME_0
timestamp 1717028433
transform 1 0 1361 0 1 -606
box -241 -384 241 384
<< labels >>
flabel metal1 1260 -2290 1460 -2180 0 FreeSans 256 0 0 0 vcont_n
port 4 nsew
flabel metal1 1260 -910 1460 -800 0 FreeSans 256 0 0 0 vcont_p
port 1 nsew
flabel metal1 1260 -2670 1460 -2560 0 FreeSans 256 0 0 0 vss
port 5 nsew
flabel metal1 1260 -320 1460 -210 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 1110 -1710 1310 -1600 0 FreeSans 256 0 0 0 in
port 3 nsew
flabel metal1 1470 -1710 1620 -1600 0 FreeSans 256 0 0 0 out
port 2 nsew
<< end >>
