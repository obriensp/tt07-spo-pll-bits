magic
tech sky130A
magscale 1 2
timestamp 1716512256
<< viali >>
rect 1508 -842 1666 -808
rect 2144 -842 2302 -808
rect 1154 -986 1312 -952
rect 1568 -986 1726 -952
rect 1056 -1552 1092 -1046
rect 2046 -1090 2204 -1056
rect 2470 -1090 2628 -1056
rect 2690 -1446 2724 -1152
<< metal1 >>
rect 1486 -280 1686 -80
rect 1812 -280 2012 -80
rect 2126 -280 2326 -80
rect 1161 -289 1219 -283
rect 1161 -606 1219 -347
rect 1554 -492 1620 -280
rect 1874 -606 1936 -280
rect 2190 -492 2256 -280
rect 2584 -332 2656 -326
rect 2584 -410 2656 -404
rect 2216 -498 2256 -492
rect 2591 -606 2649 -410
rect 1161 -664 1562 -606
rect 1608 -664 2200 -606
rect 2244 -664 2649 -606
rect 524 -808 1770 -782
rect 524 -842 1508 -808
rect 1666 -842 1770 -808
rect 524 -888 1770 -842
rect 524 -1007 618 -888
rect 524 -1194 618 -1101
rect 1044 -952 1826 -944
rect 1044 -986 1154 -952
rect 1312 -986 1568 -952
rect 1726 -986 1826 -952
rect 1044 -992 1826 -986
rect 1044 -1046 1104 -992
rect 1044 -1192 1056 -1046
rect 472 -1394 672 -1194
rect 832 -1396 1056 -1192
rect 1044 -1552 1056 -1396
rect 1092 -1192 1104 -1046
rect 1092 -1394 1210 -1192
rect 1256 -1392 1624 -1150
rect 1874 -1180 1936 -664
rect 2034 -808 2446 -790
rect 2034 -842 2144 -808
rect 2302 -842 2446 -808
rect 2034 -1050 2446 -842
rect 2822 -1016 2933 -1010
rect 1984 -1056 2730 -1050
rect 1984 -1090 2046 -1056
rect 2204 -1090 2470 -1056
rect 2628 -1090 2730 -1056
rect 1984 -1096 2730 -1090
rect 2678 -1152 2730 -1096
rect 2822 -1133 2933 -1127
rect 1674 -1356 2100 -1180
rect 2154 -1356 2522 -1182
rect 2678 -1192 2690 -1152
rect 2572 -1356 2690 -1192
rect 1092 -1552 1104 -1394
rect 1872 -1456 2158 -1396
rect 1872 -1496 1936 -1456
rect 1044 -1566 1104 -1552
rect 1200 -1702 1266 -1502
rect 1614 -1564 1936 -1496
rect 1130 -1902 1330 -1702
rect 1872 -1706 1936 -1564
rect 2516 -1704 2582 -1398
rect 2678 -1446 2690 -1356
rect 2724 -1192 2730 -1152
rect 2830 -1192 2924 -1133
rect 2724 -1356 2972 -1192
rect 2724 -1446 2730 -1356
rect 2772 -1392 2972 -1356
rect 2678 -1460 2730 -1446
rect 1814 -1906 2014 -1706
rect 2448 -1904 2648 -1704
<< via1 >>
rect 1161 -347 1219 -289
rect 2584 -404 2656 -332
rect 524 -1101 618 -1007
rect 2822 -1127 2933 -1016
<< metal2 >>
rect 1143 -356 1152 -279
rect 1229 -356 1238 -279
rect 2583 -330 2658 -321
rect 2578 -404 2583 -332
rect 2658 -404 2662 -332
rect 2583 -414 2658 -405
rect 506 -1110 515 -997
rect 628 -1110 637 -997
rect 2817 -1010 2939 -1001
rect 2816 -1127 2817 -1016
rect 2817 -1141 2939 -1132
<< via2 >>
rect 1152 -289 1229 -279
rect 1152 -347 1161 -289
rect 1161 -347 1219 -289
rect 1219 -347 1229 -289
rect 1152 -356 1229 -347
rect 2583 -332 2658 -330
rect 2583 -404 2584 -332
rect 2584 -404 2656 -332
rect 2656 -404 2658 -332
rect 2583 -405 2658 -404
rect 515 -1007 628 -997
rect 515 -1101 524 -1007
rect 524 -1101 618 -1007
rect 618 -1101 628 -1007
rect 515 -1110 628 -1101
rect 2817 -1016 2939 -1010
rect 2817 -1127 2822 -1016
rect 2822 -1127 2933 -1016
rect 2933 -1127 2939 -1016
rect 2817 -1132 2939 -1127
<< metal3 >>
rect 1147 -279 1234 -274
rect 1147 -356 1152 -279
rect 1229 -356 1234 -279
rect 1147 -361 1234 -356
rect 2578 -330 2663 -325
rect 2578 -405 2583 -330
rect 2658 -405 2663 -330
rect 2578 -410 2663 -405
rect 492 -1127 498 -980
rect 645 -1127 651 -980
rect 2809 -1001 2948 -995
rect 2809 -1146 2948 -1140
<< via3 >>
rect 498 -997 645 -980
rect 498 -1110 515 -997
rect 515 -1110 628 -997
rect 628 -1110 645 -997
rect 498 -1127 645 -1110
rect 2809 -1010 2948 -1001
rect 2809 -1132 2817 -1010
rect 2817 -1132 2939 -1010
rect 2939 -1132 2948 -1010
rect 2809 -1140 2948 -1132
<< metal4 >>
rect 498 -874 646 -470
rect 498 -979 645 -874
rect 2808 -894 2948 -496
rect 497 -980 646 -979
rect 497 -1127 498 -980
rect 645 -1127 646 -980
rect 2809 -1000 2948 -894
rect 497 -1128 646 -1127
rect 2808 -1001 2949 -1000
rect 2808 -1140 2809 -1001
rect 2948 -1140 2949 -1001
rect 2808 -1141 2949 -1140
use sky130_fd_pr__nfet_01v8_64Z3AY  sky130_fd_pr__nfet_01v8_64Z3AY_0
timestamp 1716512256
transform 1 0 2223 0 1 -599
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_LGAKDL  sky130_fd_pr__pfet_01v8_LGAKDL_0
timestamp 1716512256
transform 1 0 1647 0 1 -1300
box -211 -384 211 384
use sky130_fd_pr__cap_mim_m3_1_B4ULDW  XC1
timestamp 1716512256
transform 0 1 890 1 0 -494
box -396 -460 396 460
use sky130_fd_pr__cap_mim_m3_1_BEWQ6U  XC2
timestamp 1716512256
transform 0 1 2712 1 0 -522
box -396 -250 396 250
use sky130_fd_pr__pfet_01v8_LGAKDL  XM1
timestamp 1716512256
transform 1 0 1233 0 1 -1300
box -211 -384 211 384
use sky130_fd_pr__nfet_01v8_64QSBY  XM3
timestamp 1716512256
transform 1 0 2125 0 1 -1299
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64QSBY  XM4
timestamp 1716512256
transform 1 0 2549 0 1 -1299
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64Z3AY  XM5
timestamp 1716512256
transform 1 0 1587 0 1 -599
box -211 -279 211 279
<< labels >>
flabel metal1 832 -1392 1032 -1192 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 1814 -1906 2014 -1706 0 FreeSans 256 0 0 0 in
port 5 nsew
flabel metal1 1130 -1902 1330 -1702 0 FreeSans 256 0 0 0 vcont_p
port 1 nsew
flabel metal1 2448 -1904 2648 -1704 0 FreeSans 256 0 0 0 vcont_n
port 6 nsew
flabel metal1 1812 -280 2012 -80 0 FreeSans 256 0 0 0 out
port 4 nsew
flabel metal1 1486 -280 1686 -80 0 FreeSans 256 0 0 0 s0
port 2 nsew
flabel metal1 2126 -280 2326 -80 0 FreeSans 256 0 0 0 s1
port 3 nsew
flabel metal1 2772 -1392 2972 -1192 0 FreeSans 256 0 0 0 vss
port 7 nsew
flabel metal1 472 -1394 672 -1194 0 FreeSans 256 0 0 0 vss
port 7 nsew
<< end >>
