magic
tech sky130A
magscale 1 2
timestamp 1716512256
<< metal3 >>
rect -396 222 396 250
rect -396 -222 312 222
rect 376 -222 396 222
rect -396 -250 396 -222
<< via3 >>
rect 312 -222 376 222
<< mimcap >>
rect -356 170 64 210
rect -356 -170 -316 170
rect 24 -170 64 170
rect -356 -210 64 -170
<< mimcapcontact >>
rect -316 -170 24 170
<< metal4 >>
rect 296 222 392 238
rect -317 170 25 171
rect -317 -170 -316 170
rect 24 -170 25 170
rect -317 -171 25 -170
rect 296 -222 312 222
rect 376 -222 392 222
rect 296 -238 392 -222
<< properties >>
string FIXED_BBOX -396 -250 104 250
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.1 l 2.1 val 10.416 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
