magic
tech sky130A
magscale 1 2
timestamp 1717194565
<< error_p >>
rect -29 -207 29 -201
rect -29 -241 -17 -207
rect -29 -247 29 -241
<< pwell >>
rect -226 -379 226 379
<< nmoslvt >>
rect -30 -169 30 231
<< ndiff >>
rect -88 219 -30 231
rect -88 -157 -76 219
rect -42 -157 -30 219
rect -88 -169 -30 -157
rect 30 219 88 231
rect 30 -157 42 219
rect 76 -157 88 219
rect 30 -169 88 -157
<< ndiffc >>
rect -76 -157 -42 219
rect 42 -157 76 219
<< psubdiff >>
rect -190 309 -94 343
rect 94 309 190 343
rect -190 247 -156 309
rect 156 247 190 309
rect -190 -309 -156 -247
rect 156 -309 190 -247
rect -190 -343 -94 -309
rect 94 -343 190 -309
<< psubdiffcont >>
rect -94 309 94 343
rect -190 -247 -156 247
rect 156 -247 190 247
rect -94 -343 94 -309
<< poly >>
rect -30 231 30 257
rect -30 -191 30 -169
rect -33 -207 33 -191
rect -33 -241 -17 -207
rect 17 -241 33 -207
rect -33 -257 33 -241
<< polycont >>
rect -17 -241 17 -207
<< locali >>
rect -190 309 -94 343
rect 94 309 190 343
rect -190 247 -156 309
rect 156 247 190 309
rect -76 219 -42 235
rect -76 -173 -42 -157
rect 42 219 76 235
rect 42 -173 76 -157
rect -33 -241 -17 -207
rect 17 -241 33 -207
rect -190 -309 -156 -247
rect 156 -309 190 -247
rect -190 -343 -94 -309
rect 94 -343 190 -309
<< viali >>
rect -76 -157 -42 219
rect 42 -157 76 219
rect -17 -241 17 -207
<< metal1 >>
rect -82 219 -36 231
rect -82 -157 -76 219
rect -42 -157 -36 219
rect -82 -169 -36 -157
rect 36 219 82 231
rect 36 -157 42 219
rect 76 -157 82 219
rect 36 -169 82 -157
rect -29 -207 29 -201
rect -29 -241 -17 -207
rect 17 -241 29 -207
rect -29 -247 29 -241
<< properties >>
string FIXED_BBOX -173 -326 173 326
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
